VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

# High density, single height
SITE obssite
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.36 BY 6.12 ;
END obssite

#--------EOF---------

MACRO AN2D1
  CLASS CORE ;
  FOREIGN AN2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 3.435 1.090 3.605 4.220 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 5.400 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.400 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 5.400 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 5.400 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 5.580 6.445 ;
      LAYER pwell ;
        RECT 3.245 1.625 4.875 1.690 ;
        RECT 0.005 0.730 4.875 1.625 ;
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 1.275 3.230 1.445 4.220 ;
        RECT 1.275 3.060 2.605 3.230 ;
        RECT 2.355 1.090 2.525 3.060 ;
        RECT 2.275 0.920 2.605 1.090 ;
  END
END AN2D1

#--------EOF---------

MACRO AN2D1_1
  CLASS CORE ;
  FOREIGN AN2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 3.435 1.090 3.605 4.220 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 1.735 1.980 2.065 2.150 ;
        RECT 1.815 1.330 1.985 1.980 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.320 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 4.320 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 4.320 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 4.500 6.445 ;
      LAYER pwell ;
        RECT 2.165 1.625 3.795 1.690 ;
        RECT 0.005 0.730 3.795 1.625 ;
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 1.275 3.230 1.445 4.220 ;
        RECT 1.275 3.060 3.145 3.230 ;
        RECT 1.275 2.690 1.445 3.060 ;
        RECT 1.275 2.520 3.145 2.690 ;
        RECT 1.275 1.090 1.445 2.520 ;
        RECT 0.115 0.920 1.445 1.090 ;
  END
END AN2D1_1

#--------EOF---------

MACRO AN2D1_2
  CLASS CORE ;
  FOREIGN AN2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 3.435 1.090 3.605 4.220 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 5.400 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.400 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 5.400 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 5.400 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 5.580 6.445 ;
      LAYER pwell ;
        RECT 3.245 1.625 4.875 1.690 ;
        RECT 0.005 0.730 4.875 1.625 ;
      LAYER li1 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 2.275 4.220 2.605 4.390 ;
        RECT 0.195 3.230 0.365 4.220 ;
        RECT 2.355 3.230 2.525 4.220 ;
        RECT 0.195 3.060 2.605 3.230 ;
        RECT 2.355 1.090 2.525 3.060 ;
        RECT 2.275 0.920 2.605 1.090 ;
  END
END AN2D1_2

#--------EOF---------

MACRO AN2D1_3
  CLASS CORE ;
  FOREIGN AN2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 3.435 1.090 3.605 4.220 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 5.400 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.400 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 5.400 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 5.400 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 5.580 6.445 ;
      LAYER pwell ;
        RECT 3.245 1.625 4.875 1.690 ;
        RECT 0.005 0.730 4.875 1.625 ;
      LAYER li1 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 2.275 4.220 2.605 4.390 ;
        RECT 0.195 3.230 0.365 4.220 ;
        RECT 2.355 3.230 2.525 4.220 ;
        RECT 0.195 3.060 2.605 3.230 ;
        RECT 0.195 1.090 0.365 3.060 ;
        RECT 0.115 0.920 0.445 1.090 ;
  END
END AN2D1_3

#--------EOF---------

MACRO AO21D1
  CLASS CORE ;
  FOREIGN AO21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 4.435 4.220 4.765 4.390 ;
        RECT 4.515 1.090 4.685 4.220 ;
        RECT 4.435 0.920 4.765 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 0.000 -0.085 6.480 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.480 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 6.480 6.205 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 6.480 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 6.660 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 5.955 1.690 ;
      LAYER li1 ;
        RECT 0.115 4.220 2.605 4.390 ;
        RECT 1.275 3.230 1.445 4.220 ;
        RECT 0.195 3.060 4.225 3.230 ;
        RECT 0.195 1.090 0.365 3.060 ;
        RECT 3.435 1.090 3.605 3.060 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 3.435 0.440 3.605 0.920 ;
        RECT 3.435 0.270 5.305 0.440 ;
  END
END AO21D1

#--------EOF---------

MACRO AO21D1_1
  CLASS CORE ;
  FOREIGN AO21D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 3.975 2.150 4.145 2.690 ;
        RECT 3.895 1.980 4.225 2.150 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 5.515 4.220 5.845 4.390 ;
        RECT 5.595 1.090 5.765 4.220 ;
        RECT 5.515 0.920 5.845 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 6.480 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.480 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 6.480 6.205 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 6.480 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 6.660 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 5.955 1.690 ;
      LAYER li1 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 1.195 4.220 3.685 4.390 ;
        RECT 0.195 3.230 0.365 4.220 ;
        RECT 2.355 3.230 2.525 4.220 ;
        RECT 0.195 3.060 2.525 3.230 ;
        RECT 2.355 1.090 2.525 3.060 ;
        RECT 2.275 0.920 3.685 1.090 ;
        RECT 2.355 0.440 2.525 0.920 ;
        RECT 2.275 0.270 2.605 0.440 ;
  END
END AO21D1_1

#--------EOF---------

MACRO AO21D1_2
  CLASS CORE ;
  FOREIGN AO21D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.195 2.150 0.365 2.690 ;
        RECT 0.115 1.980 0.445 2.150 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 4.435 4.220 4.765 4.390 ;
        RECT 4.515 1.090 4.685 4.220 ;
        RECT 4.435 0.920 4.765 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 0.000 -0.085 6.480 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.480 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 6.480 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 6.480 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 6.660 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 5.955 1.690 ;
      LAYER li1 ;
        RECT 0.735 4.690 2.605 4.860 ;
        RECT 0.735 1.090 0.905 4.690 ;
        RECT 1.195 4.220 3.685 4.390 ;
        RECT 0.735 0.920 1.525 1.090 ;
        RECT 1.275 0.440 1.445 0.920 ;
        RECT 1.195 0.270 1.525 0.440 ;
  END
END AO21D1_2

#--------EOF---------

MACRO AO21D1_3
  CLASS CORE ;
  FOREIGN AO21D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 4.435 4.220 4.765 4.390 ;
        RECT 4.515 1.090 4.685 4.220 ;
        RECT 4.435 0.920 4.765 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 0.000 -0.085 6.480 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.480 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 6.480 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 6.480 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 6.660 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 5.955 1.690 ;
      LAYER li1 ;
        RECT 1.195 4.220 3.685 4.390 ;
        RECT 2.355 3.230 2.525 4.220 ;
        RECT 2.355 3.060 3.605 3.230 ;
        RECT 3.435 1.090 3.605 3.060 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 0.195 0.440 0.365 0.920 ;
        RECT 3.435 0.440 3.605 0.920 ;
        RECT 0.115 0.270 0.445 0.440 ;
        RECT 3.435 0.270 5.305 0.440 ;
  END
END AO21D1_3

#--------EOF---------

MACRO AOI21D1
  CLASS CORE ;
  FOREIGN AOI21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.368000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 4.220 2.605 4.390 ;
        RECT 1.275 3.230 1.445 4.220 ;
        RECT 1.275 3.060 2.525 3.230 ;
        RECT 2.355 1.090 2.525 3.060 ;
        RECT 2.275 0.920 2.605 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.320 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 4.320 6.205 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 3.355 5.030 3.685 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 4.320 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 4.500 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 3.795 1.690 ;
  END
END AOI21D1

#--------EOF---------

MACRO AOI21D1_1
  CLASS CORE ;
  FOREIGN AOI21D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.368000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 3.685 4.390 ;
        RECT 2.355 3.230 2.525 4.220 ;
        RECT 1.275 3.060 2.525 3.230 ;
        RECT 1.275 1.090 1.445 3.060 ;
        RECT 1.195 0.920 1.525 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.320 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 4.320 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 4.320 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 4.500 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 3.795 1.690 ;
  END
END AOI21D1_1

#--------EOF---------

MACRO AOI21D1_2
  CLASS CORE ;
  FOREIGN AOI21D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.890000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 1.195 4.220 3.685 4.390 ;
        RECT 0.195 3.230 0.365 4.220 ;
        RECT 2.355 3.230 2.525 4.220 ;
        RECT 0.195 3.060 2.525 3.230 ;
        RECT 2.355 1.090 2.525 3.060 ;
        RECT 2.275 0.920 3.685 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 3.975 2.150 4.145 2.690 ;
        RECT 3.895 1.980 4.225 2.150 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 5.400 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.400 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 5.400 6.205 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 5.400 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 5.580 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 4.875 1.690 ;
  END
END AOI21D1_2

#--------EOF---------

MACRO AOI21D1_3
  CLASS CORE ;
  FOREIGN AOI21D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.890000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 1.195 4.220 3.685 4.390 ;
        RECT 0.195 3.230 0.365 4.220 ;
        RECT 2.355 3.230 2.525 4.220 ;
        RECT 0.195 3.060 2.525 3.230 ;
        RECT 0.195 2.690 0.365 3.060 ;
        RECT 0.195 2.520 3.605 2.690 ;
        RECT 0.195 1.090 0.365 2.520 ;
        RECT 3.435 1.090 3.605 2.520 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.980 0.985 2.150 ;
        RECT 0.735 1.330 0.905 1.980 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.735 1.980 2.065 2.150 ;
        RECT 1.815 1.330 1.985 1.980 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 3.975 2.150 4.145 2.690 ;
        RECT 3.895 1.980 4.225 2.150 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 5.400 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.400 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 5.400 6.205 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 5.400 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 5.580 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 4.875 1.690 ;
  END
END AOI21D1_3

#--------EOF---------

MACRO BUFFD1
  CLASS CORE ;
  FOREIGN BUFFD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 0.195 1.090 0.365 4.220 ;
        RECT 0.115 0.920 0.445 1.090 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.145500 ;
    PORT
      LAYER li1 ;
        RECT 2.355 2.690 2.525 3.230 ;
        RECT 2.275 2.520 2.605 2.690 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 0.000 -0.085 3.240 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.240 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 3.240 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 3.240 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 3.420 6.445 ;
      LAYER pwell ;
        RECT 0.005 1.410 1.635 1.690 ;
        RECT 0.005 0.730 2.715 1.410 ;
      LAYER li1 ;
        RECT 1.815 5.030 2.605 5.200 ;
        RECT 1.815 3.230 1.985 5.030 ;
        RECT 1.735 3.060 2.065 3.230 ;
        RECT 0.655 1.980 2.525 2.150 ;
        RECT 2.355 1.090 2.525 1.980 ;
        RECT 2.275 0.920 2.605 1.090 ;
  END
END BUFFD1

#--------EOF---------

MACRO BUFFD1_1
  CLASS CORE ;
  FOREIGN BUFFD1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 4.220 2.605 4.390 ;
        RECT 2.355 1.090 2.525 4.220 ;
        RECT 2.275 0.920 2.605 1.090 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.145500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 4.220 0.985 4.390 ;
        RECT 0.735 0.440 0.905 4.220 ;
        RECT 0.655 0.270 0.985 0.440 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 0.000 -0.085 3.240 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.240 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 3.240 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 3.240 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 3.420 6.445 ;
      LAYER pwell ;
        RECT 1.085 1.410 2.715 1.690 ;
        RECT 0.005 0.730 2.715 1.410 ;
      LAYER li1 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 0.195 3.230 0.365 5.030 ;
        RECT 0.115 3.060 0.445 3.230 ;
        RECT 0.115 1.980 0.445 2.150 ;
        RECT 0.195 1.090 0.365 1.980 ;
        RECT 0.115 0.920 0.445 1.090 ;
  END
END BUFFD1_1

#--------EOF---------

MACRO DFCNQD1
  CLASS CORE ;
  FOREIGN DFCNQD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.184500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END d
  PIN cdn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.379500 ;
    PORT
      LAYER li1 ;
        RECT 4.515 0.270 5.305 0.440 ;
    END
  END cdn
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.145500 ;
    PORT
      LAYER li1 ;
        RECT 6.055 1.980 6.845 2.150 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 17.395 4.220 17.725 4.390 ;
        RECT 17.475 1.090 17.645 4.220 ;
        RECT 17.395 0.920 17.725 1.090 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 8.755 0.920 9.085 1.090 ;
        RECT 13.075 0.920 13.405 1.090 ;
        RECT 18.475 0.920 18.805 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 8.835 0.085 9.005 0.920 ;
        RECT 13.155 0.085 13.325 0.920 ;
        RECT 18.555 0.085 18.725 0.920 ;
        RECT 0.000 -0.085 19.440 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
        RECT 10.895 -0.085 11.065 0.085 ;
        RECT 11.255 -0.085 11.425 0.085 ;
        RECT 11.615 -0.085 11.785 0.085 ;
        RECT 11.975 -0.085 12.145 0.085 ;
        RECT 12.335 -0.085 12.505 0.085 ;
        RECT 12.695 -0.085 12.865 0.085 ;
        RECT 13.055 -0.085 13.225 0.085 ;
        RECT 13.415 -0.085 13.585 0.085 ;
        RECT 13.775 -0.085 13.945 0.085 ;
        RECT 14.135 -0.085 14.305 0.085 ;
        RECT 14.495 -0.085 14.665 0.085 ;
        RECT 14.855 -0.085 15.025 0.085 ;
        RECT 15.215 -0.085 15.385 0.085 ;
        RECT 15.575 -0.085 15.745 0.085 ;
        RECT 15.935 -0.085 16.105 0.085 ;
        RECT 16.295 -0.085 16.465 0.085 ;
        RECT 16.655 -0.085 16.825 0.085 ;
        RECT 17.015 -0.085 17.185 0.085 ;
        RECT 17.375 -0.085 17.545 0.085 ;
        RECT 17.735 -0.085 17.905 0.085 ;
        RECT 18.095 -0.085 18.265 0.085 ;
        RECT 18.455 -0.085 18.625 0.085 ;
        RECT 18.815 -0.085 18.985 0.085 ;
        RECT 19.175 -0.085 19.345 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 19.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 19.440 6.205 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 8.835 5.200 9.005 6.035 ;
        RECT 13.155 5.200 13.325 6.035 ;
        RECT 16.395 5.200 16.565 6.035 ;
        RECT 18.555 5.200 18.725 6.035 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 8.755 5.030 9.085 5.200 ;
        RECT 13.075 5.030 13.405 5.200 ;
        RECT 16.315 5.030 16.645 5.200 ;
        RECT 18.475 5.030 18.805 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
        RECT 10.895 6.035 11.065 6.205 ;
        RECT 11.255 6.035 11.425 6.205 ;
        RECT 11.615 6.035 11.785 6.205 ;
        RECT 11.975 6.035 12.145 6.205 ;
        RECT 12.335 6.035 12.505 6.205 ;
        RECT 12.695 6.035 12.865 6.205 ;
        RECT 13.055 6.035 13.225 6.205 ;
        RECT 13.415 6.035 13.585 6.205 ;
        RECT 13.775 6.035 13.945 6.205 ;
        RECT 14.135 6.035 14.305 6.205 ;
        RECT 14.495 6.035 14.665 6.205 ;
        RECT 14.855 6.035 15.025 6.205 ;
        RECT 15.215 6.035 15.385 6.205 ;
        RECT 15.575 6.035 15.745 6.205 ;
        RECT 15.935 6.035 16.105 6.205 ;
        RECT 16.295 6.035 16.465 6.205 ;
        RECT 16.655 6.035 16.825 6.205 ;
        RECT 17.015 6.035 17.185 6.205 ;
        RECT 17.375 6.035 17.545 6.205 ;
        RECT 17.735 6.035 17.905 6.205 ;
        RECT 18.095 6.035 18.265 6.205 ;
        RECT 18.455 6.035 18.625 6.205 ;
        RECT 18.815 6.035 18.985 6.205 ;
        RECT 19.175 6.035 19.345 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 19.440 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 19.620 6.445 ;
      LAYER pwell ;
        RECT 7.565 1.480 9.195 1.690 ;
        RECT 7.565 1.410 11.355 1.480 ;
        RECT 15.125 1.410 18.915 1.690 ;
        RECT 0.005 0.730 18.915 1.410 ;
      LAYER li1 ;
        RECT 0.115 5.030 3.065 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
        RECT 14.155 5.030 14.485 5.200 ;
        RECT 2.895 4.860 3.065 5.030 ;
        RECT 4.515 4.860 4.685 5.030 ;
        RECT 1.195 4.690 1.525 4.860 ;
        RECT 2.895 4.690 4.685 4.860 ;
        RECT 10.915 4.690 11.705 4.860 ;
        RECT 1.275 4.390 1.445 4.690 ;
        RECT 1.275 4.220 2.525 4.390 ;
        RECT 2.355 1.090 2.525 4.220 ;
        RECT 11.535 3.230 11.705 4.690 ;
        RECT 14.235 4.390 14.405 5.030 ;
        RECT 11.995 4.220 14.405 4.390 ;
        RECT 11.455 3.060 11.785 3.230 ;
        RECT 14.235 2.690 14.405 4.220 ;
        RECT 3.975 2.520 10.165 2.690 ;
        RECT 14.155 2.520 14.485 2.690 ;
        RECT 3.975 2.150 4.145 2.520 ;
        RECT 2.815 1.980 4.145 2.150 ;
        RECT 7.755 1.980 9.625 2.150 ;
        RECT 7.755 1.500 7.925 1.980 ;
        RECT 5.055 1.330 7.925 1.500 ;
        RECT 8.295 1.330 16.565 1.500 ;
        RECT 5.055 1.090 5.225 1.330 ;
        RECT 8.295 1.090 8.465 1.330 ;
        RECT 16.395 1.090 16.565 1.330 ;
        RECT 2.275 0.920 5.225 1.090 ;
        RECT 7.675 0.920 8.465 1.090 ;
        RECT 10.915 0.920 12.785 1.090 ;
        RECT 14.155 0.920 15.025 1.090 ;
        RECT 16.315 0.920 16.645 1.090 ;
        RECT 12.615 0.440 12.785 0.920 ;
        RECT 12.535 0.270 12.865 0.440 ;
  END
END DFCNQD1

#--------EOF---------

MACRO DFCNQD1_1
  CLASS CORE ;
  FOREIGN DFCNQD1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.184500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END d
  PIN cdn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.379500 ;
    PORT
      LAYER li1 ;
        RECT 4.515 0.270 5.305 0.440 ;
    END
  END cdn
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.145500 ;
    PORT
      LAYER li1 ;
        RECT 6.055 1.980 6.845 2.150 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 14.155 4.220 14.485 4.390 ;
        RECT 14.235 1.090 14.405 4.220 ;
        RECT 14.155 0.920 14.485 1.090 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 8.755 0.920 9.085 1.090 ;
        RECT 13.075 0.920 13.405 1.090 ;
        RECT 18.475 0.920 18.805 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 8.835 0.085 9.005 0.920 ;
        RECT 13.155 0.085 13.325 0.920 ;
        RECT 18.555 0.085 18.725 0.920 ;
        RECT 0.000 -0.085 19.440 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
        RECT 10.895 -0.085 11.065 0.085 ;
        RECT 11.255 -0.085 11.425 0.085 ;
        RECT 11.615 -0.085 11.785 0.085 ;
        RECT 11.975 -0.085 12.145 0.085 ;
        RECT 12.335 -0.085 12.505 0.085 ;
        RECT 12.695 -0.085 12.865 0.085 ;
        RECT 13.055 -0.085 13.225 0.085 ;
        RECT 13.415 -0.085 13.585 0.085 ;
        RECT 13.775 -0.085 13.945 0.085 ;
        RECT 14.135 -0.085 14.305 0.085 ;
        RECT 14.495 -0.085 14.665 0.085 ;
        RECT 14.855 -0.085 15.025 0.085 ;
        RECT 15.215 -0.085 15.385 0.085 ;
        RECT 15.575 -0.085 15.745 0.085 ;
        RECT 15.935 -0.085 16.105 0.085 ;
        RECT 16.295 -0.085 16.465 0.085 ;
        RECT 16.655 -0.085 16.825 0.085 ;
        RECT 17.015 -0.085 17.185 0.085 ;
        RECT 17.375 -0.085 17.545 0.085 ;
        RECT 17.735 -0.085 17.905 0.085 ;
        RECT 18.095 -0.085 18.265 0.085 ;
        RECT 18.455 -0.085 18.625 0.085 ;
        RECT 18.815 -0.085 18.985 0.085 ;
        RECT 19.175 -0.085 19.345 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 19.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 19.440 6.205 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 8.835 5.200 9.005 6.035 ;
        RECT 13.155 5.200 13.325 6.035 ;
        RECT 16.395 5.200 16.565 6.035 ;
        RECT 18.555 5.200 18.725 6.035 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 8.755 5.030 9.085 5.200 ;
        RECT 13.075 5.030 13.405 5.200 ;
        RECT 16.315 5.030 16.645 5.200 ;
        RECT 18.475 5.030 18.805 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
        RECT 10.895 6.035 11.065 6.205 ;
        RECT 11.255 6.035 11.425 6.205 ;
        RECT 11.615 6.035 11.785 6.205 ;
        RECT 11.975 6.035 12.145 6.205 ;
        RECT 12.335 6.035 12.505 6.205 ;
        RECT 12.695 6.035 12.865 6.205 ;
        RECT 13.055 6.035 13.225 6.205 ;
        RECT 13.415 6.035 13.585 6.205 ;
        RECT 13.775 6.035 13.945 6.205 ;
        RECT 14.135 6.035 14.305 6.205 ;
        RECT 14.495 6.035 14.665 6.205 ;
        RECT 14.855 6.035 15.025 6.205 ;
        RECT 15.215 6.035 15.385 6.205 ;
        RECT 15.575 6.035 15.745 6.205 ;
        RECT 15.935 6.035 16.105 6.205 ;
        RECT 16.295 6.035 16.465 6.205 ;
        RECT 16.655 6.035 16.825 6.205 ;
        RECT 17.015 6.035 17.185 6.205 ;
        RECT 17.375 6.035 17.545 6.205 ;
        RECT 17.735 6.035 17.905 6.205 ;
        RECT 18.095 6.035 18.265 6.205 ;
        RECT 18.455 6.035 18.625 6.205 ;
        RECT 18.815 6.035 18.985 6.205 ;
        RECT 19.175 6.035 19.345 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 19.440 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 19.620 6.445 ;
      LAYER pwell ;
        RECT 7.565 1.480 9.195 1.690 ;
        RECT 7.565 1.410 11.355 1.480 ;
        RECT 12.965 1.410 16.755 1.690 ;
        RECT 0.005 0.730 18.915 1.410 ;
      LAYER li1 ;
        RECT 11.455 5.680 11.785 5.850 ;
        RECT 11.535 5.200 11.705 5.680 ;
        RECT 0.115 5.030 3.065 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
        RECT 9.915 5.030 11.705 5.200 ;
        RECT 16.935 5.030 17.725 5.200 ;
        RECT 2.895 4.860 3.065 5.030 ;
        RECT 4.515 4.860 4.685 5.030 ;
        RECT 1.195 4.690 1.525 4.860 ;
        RECT 2.895 4.690 4.685 4.860 ;
        RECT 1.275 4.390 1.445 4.690 ;
        RECT 1.275 4.220 2.525 4.390 ;
        RECT 2.355 1.090 2.525 4.220 ;
        RECT 9.915 2.690 10.085 5.030 ;
        RECT 10.915 4.690 11.705 4.860 ;
        RECT 11.535 3.230 11.705 4.690 ;
        RECT 11.455 3.060 11.785 3.230 ;
        RECT 3.975 2.520 10.165 2.690 ;
        RECT 3.975 2.150 4.145 2.520 ;
        RECT 16.935 2.150 17.105 5.030 ;
        RECT 2.815 1.980 4.145 2.150 ;
        RECT 7.755 1.980 9.625 2.150 ;
        RECT 15.235 1.980 17.105 2.150 ;
        RECT 7.755 1.500 7.925 1.980 ;
        RECT 5.055 1.330 7.925 1.500 ;
        RECT 8.295 1.330 13.865 1.500 ;
        RECT 5.055 1.090 5.225 1.330 ;
        RECT 8.295 1.090 8.465 1.330 ;
        RECT 2.275 0.920 5.225 1.090 ;
        RECT 7.675 0.920 8.465 1.090 ;
        RECT 10.915 0.920 12.785 1.090 ;
        RECT 12.615 0.440 12.785 0.920 ;
        RECT 13.695 0.440 13.865 1.330 ;
        RECT 16.935 1.090 17.105 1.980 ;
        RECT 16.315 0.920 16.645 1.090 ;
        RECT 16.935 0.920 17.725 1.090 ;
        RECT 16.395 0.440 16.565 0.920 ;
        RECT 12.535 0.270 12.865 0.440 ;
        RECT 13.695 0.270 16.565 0.440 ;
  END
END DFCNQD1_1

#--------EOF---------

MACRO DFCNQD1_2
  CLASS CORE ;
  FOREIGN DFCNQD1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.184500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END d
  PIN cdn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.379500 ;
    PORT
      LAYER li1 ;
        RECT 4.515 0.270 5.305 0.440 ;
    END
  END cdn
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.145500 ;
    PORT
      LAYER li1 ;
        RECT 6.055 1.980 6.845 2.150 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 17.395 4.220 17.725 4.390 ;
        RECT 17.475 1.090 17.645 4.220 ;
        RECT 17.395 0.920 17.725 1.090 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 8.755 0.920 9.085 1.090 ;
        RECT 13.075 0.920 13.405 1.090 ;
        RECT 18.475 0.920 18.805 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 8.835 0.085 9.005 0.920 ;
        RECT 13.155 0.085 13.325 0.920 ;
        RECT 18.555 0.085 18.725 0.920 ;
        RECT 0.000 -0.085 19.440 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
        RECT 10.895 -0.085 11.065 0.085 ;
        RECT 11.255 -0.085 11.425 0.085 ;
        RECT 11.615 -0.085 11.785 0.085 ;
        RECT 11.975 -0.085 12.145 0.085 ;
        RECT 12.335 -0.085 12.505 0.085 ;
        RECT 12.695 -0.085 12.865 0.085 ;
        RECT 13.055 -0.085 13.225 0.085 ;
        RECT 13.415 -0.085 13.585 0.085 ;
        RECT 13.775 -0.085 13.945 0.085 ;
        RECT 14.135 -0.085 14.305 0.085 ;
        RECT 14.495 -0.085 14.665 0.085 ;
        RECT 14.855 -0.085 15.025 0.085 ;
        RECT 15.215 -0.085 15.385 0.085 ;
        RECT 15.575 -0.085 15.745 0.085 ;
        RECT 15.935 -0.085 16.105 0.085 ;
        RECT 16.295 -0.085 16.465 0.085 ;
        RECT 16.655 -0.085 16.825 0.085 ;
        RECT 17.015 -0.085 17.185 0.085 ;
        RECT 17.375 -0.085 17.545 0.085 ;
        RECT 17.735 -0.085 17.905 0.085 ;
        RECT 18.095 -0.085 18.265 0.085 ;
        RECT 18.455 -0.085 18.625 0.085 ;
        RECT 18.815 -0.085 18.985 0.085 ;
        RECT 19.175 -0.085 19.345 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 19.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 19.440 6.205 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 8.835 5.200 9.005 6.035 ;
        RECT 13.155 5.200 13.325 6.035 ;
        RECT 16.395 5.200 16.565 6.035 ;
        RECT 18.555 5.200 18.725 6.035 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 8.755 5.030 9.085 5.200 ;
        RECT 13.075 5.030 13.405 5.200 ;
        RECT 16.315 5.030 16.645 5.200 ;
        RECT 18.475 5.030 18.805 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
        RECT 10.895 6.035 11.065 6.205 ;
        RECT 11.255 6.035 11.425 6.205 ;
        RECT 11.615 6.035 11.785 6.205 ;
        RECT 11.975 6.035 12.145 6.205 ;
        RECT 12.335 6.035 12.505 6.205 ;
        RECT 12.695 6.035 12.865 6.205 ;
        RECT 13.055 6.035 13.225 6.205 ;
        RECT 13.415 6.035 13.585 6.205 ;
        RECT 13.775 6.035 13.945 6.205 ;
        RECT 14.135 6.035 14.305 6.205 ;
        RECT 14.495 6.035 14.665 6.205 ;
        RECT 14.855 6.035 15.025 6.205 ;
        RECT 15.215 6.035 15.385 6.205 ;
        RECT 15.575 6.035 15.745 6.205 ;
        RECT 15.935 6.035 16.105 6.205 ;
        RECT 16.295 6.035 16.465 6.205 ;
        RECT 16.655 6.035 16.825 6.205 ;
        RECT 17.015 6.035 17.185 6.205 ;
        RECT 17.375 6.035 17.545 6.205 ;
        RECT 17.735 6.035 17.905 6.205 ;
        RECT 18.095 6.035 18.265 6.205 ;
        RECT 18.455 6.035 18.625 6.205 ;
        RECT 18.815 6.035 18.985 6.205 ;
        RECT 19.175 6.035 19.345 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 19.440 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 19.620 6.445 ;
      LAYER pwell ;
        RECT 7.565 1.410 9.195 1.690 ;
        RECT 10.805 1.420 12.435 1.480 ;
        RECT 10.805 1.410 13.515 1.420 ;
        RECT 15.125 1.410 18.915 1.690 ;
        RECT 0.005 0.730 18.915 1.410 ;
      LAYER li1 ;
        RECT 0.115 5.030 3.065 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
        RECT 14.155 5.030 14.485 5.200 ;
        RECT 2.895 4.860 3.065 5.030 ;
        RECT 4.515 4.860 4.685 5.030 ;
        RECT 1.195 4.690 1.525 4.860 ;
        RECT 2.895 4.690 4.685 4.860 ;
        RECT 10.915 4.690 11.705 4.860 ;
        RECT 1.275 4.390 1.445 4.690 ;
        RECT 1.275 4.220 2.525 4.390 ;
        RECT 2.355 1.090 2.525 4.220 ;
        RECT 11.535 3.230 11.705 4.690 ;
        RECT 11.535 3.060 13.405 3.230 ;
        RECT 14.235 2.690 14.405 5.030 ;
        RECT 3.975 2.520 9.085 2.690 ;
        RECT 11.995 2.520 14.945 2.690 ;
        RECT 3.975 2.150 4.145 2.520 ;
        RECT 14.775 2.150 14.945 2.520 ;
        RECT 2.815 1.980 4.145 2.150 ;
        RECT 7.755 1.980 12.865 2.150 ;
        RECT 14.695 1.980 15.025 2.150 ;
        RECT 7.755 1.500 7.925 1.980 ;
        RECT 5.055 1.330 7.925 1.500 ;
        RECT 8.295 1.330 16.565 1.500 ;
        RECT 5.055 1.090 5.225 1.330 ;
        RECT 8.295 1.090 8.465 1.330 ;
        RECT 16.395 1.090 16.565 1.330 ;
        RECT 2.275 0.920 5.225 1.090 ;
        RECT 7.675 0.920 8.465 1.090 ;
        RECT 10.915 0.920 12.785 1.090 ;
        RECT 14.155 0.920 15.025 1.090 ;
        RECT 16.315 0.920 16.645 1.090 ;
        RECT 12.615 0.440 12.785 0.920 ;
        RECT 12.535 0.270 12.865 0.440 ;
  END
END DFCNQD1_2

#--------EOF---------

MACRO DFCNQD1_3
  CLASS CORE ;
  FOREIGN DFCNQD1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.184500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END d
  PIN cdn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.379500 ;
    PORT
      LAYER li1 ;
        RECT 4.515 0.270 5.305 0.440 ;
    END
  END cdn
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.145500 ;
    PORT
      LAYER li1 ;
        RECT 6.055 1.980 6.845 2.150 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 14.155 4.220 14.485 4.390 ;
        RECT 14.235 1.090 14.405 4.220 ;
        RECT 14.155 0.920 14.485 1.090 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 8.755 0.920 9.085 1.090 ;
        RECT 13.075 0.920 13.405 1.090 ;
        RECT 18.475 0.920 18.805 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 8.835 0.085 9.005 0.920 ;
        RECT 13.155 0.085 13.325 0.920 ;
        RECT 18.555 0.085 18.725 0.920 ;
        RECT 0.000 -0.085 19.440 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
        RECT 10.895 -0.085 11.065 0.085 ;
        RECT 11.255 -0.085 11.425 0.085 ;
        RECT 11.615 -0.085 11.785 0.085 ;
        RECT 11.975 -0.085 12.145 0.085 ;
        RECT 12.335 -0.085 12.505 0.085 ;
        RECT 12.695 -0.085 12.865 0.085 ;
        RECT 13.055 -0.085 13.225 0.085 ;
        RECT 13.415 -0.085 13.585 0.085 ;
        RECT 13.775 -0.085 13.945 0.085 ;
        RECT 14.135 -0.085 14.305 0.085 ;
        RECT 14.495 -0.085 14.665 0.085 ;
        RECT 14.855 -0.085 15.025 0.085 ;
        RECT 15.215 -0.085 15.385 0.085 ;
        RECT 15.575 -0.085 15.745 0.085 ;
        RECT 15.935 -0.085 16.105 0.085 ;
        RECT 16.295 -0.085 16.465 0.085 ;
        RECT 16.655 -0.085 16.825 0.085 ;
        RECT 17.015 -0.085 17.185 0.085 ;
        RECT 17.375 -0.085 17.545 0.085 ;
        RECT 17.735 -0.085 17.905 0.085 ;
        RECT 18.095 -0.085 18.265 0.085 ;
        RECT 18.455 -0.085 18.625 0.085 ;
        RECT 18.815 -0.085 18.985 0.085 ;
        RECT 19.175 -0.085 19.345 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 19.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 19.440 6.205 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 8.835 5.200 9.005 6.035 ;
        RECT 13.155 5.200 13.325 6.035 ;
        RECT 16.395 5.200 16.565 6.035 ;
        RECT 18.555 5.200 18.725 6.035 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 8.755 5.030 9.085 5.200 ;
        RECT 13.075 5.030 13.405 5.200 ;
        RECT 16.315 5.030 16.645 5.200 ;
        RECT 18.475 5.030 18.805 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
        RECT 10.895 6.035 11.065 6.205 ;
        RECT 11.255 6.035 11.425 6.205 ;
        RECT 11.615 6.035 11.785 6.205 ;
        RECT 11.975 6.035 12.145 6.205 ;
        RECT 12.335 6.035 12.505 6.205 ;
        RECT 12.695 6.035 12.865 6.205 ;
        RECT 13.055 6.035 13.225 6.205 ;
        RECT 13.415 6.035 13.585 6.205 ;
        RECT 13.775 6.035 13.945 6.205 ;
        RECT 14.135 6.035 14.305 6.205 ;
        RECT 14.495 6.035 14.665 6.205 ;
        RECT 14.855 6.035 15.025 6.205 ;
        RECT 15.215 6.035 15.385 6.205 ;
        RECT 15.575 6.035 15.745 6.205 ;
        RECT 15.935 6.035 16.105 6.205 ;
        RECT 16.295 6.035 16.465 6.205 ;
        RECT 16.655 6.035 16.825 6.205 ;
        RECT 17.015 6.035 17.185 6.205 ;
        RECT 17.375 6.035 17.545 6.205 ;
        RECT 17.735 6.035 17.905 6.205 ;
        RECT 18.095 6.035 18.265 6.205 ;
        RECT 18.455 6.035 18.625 6.205 ;
        RECT 18.815 6.035 18.985 6.205 ;
        RECT 19.175 6.035 19.345 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 19.440 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 19.620 6.445 ;
      LAYER pwell ;
        RECT 7.565 1.410 9.195 1.690 ;
        RECT 12.965 1.480 16.755 1.690 ;
        RECT 10.805 1.410 16.755 1.480 ;
        RECT 0.005 0.730 18.915 1.410 ;
      LAYER li1 ;
        RECT 0.115 5.030 3.065 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
        RECT 16.935 5.030 17.725 5.200 ;
        RECT 2.895 4.860 3.065 5.030 ;
        RECT 4.515 4.860 4.685 5.030 ;
        RECT 1.195 4.690 1.525 4.860 ;
        RECT 2.895 4.690 4.685 4.860 ;
        RECT 10.915 4.690 11.705 4.860 ;
        RECT 1.275 4.390 1.445 4.690 ;
        RECT 1.275 4.220 2.525 4.390 ;
        RECT 2.355 1.090 2.525 4.220 ;
        RECT 11.535 3.230 11.705 4.690 ;
        RECT 11.535 3.060 13.405 3.230 ;
        RECT 16.935 2.690 17.105 5.030 ;
        RECT 3.975 2.520 9.085 2.690 ;
        RECT 11.995 2.520 13.945 2.690 ;
        RECT 15.235 2.520 17.105 2.690 ;
        RECT 3.975 2.150 4.145 2.520 ;
        RECT 2.815 1.980 4.145 2.150 ;
        RECT 7.755 1.980 12.865 2.150 ;
        RECT 7.755 1.500 7.925 1.980 ;
        RECT 5.055 1.330 7.925 1.500 ;
        RECT 8.295 1.330 13.865 1.500 ;
        RECT 5.055 1.090 5.225 1.330 ;
        RECT 8.295 1.090 8.465 1.330 ;
        RECT 2.275 0.920 5.225 1.090 ;
        RECT 7.675 0.920 8.465 1.090 ;
        RECT 10.915 0.920 12.785 1.090 ;
        RECT 12.615 0.440 12.785 0.920 ;
        RECT 13.695 0.440 13.865 1.330 ;
        RECT 16.935 1.090 17.105 2.520 ;
        RECT 16.315 0.920 16.645 1.090 ;
        RECT 16.935 0.920 17.725 1.090 ;
        RECT 16.395 0.440 16.565 0.920 ;
        RECT 12.535 0.270 12.865 0.440 ;
        RECT 13.695 0.270 16.565 0.440 ;
  END
END DFCNQD1_3

#--------EOF---------

MACRO DFQD1
  CLASS CORE ;
  FOREIGN DFQD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.280 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.166500 ;
    PORT
      LAYER li1 ;
        RECT 2.815 1.980 3.145 2.150 ;
        RECT 2.895 1.330 3.065 1.980 ;
    END
  END d
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 15.235 4.220 15.565 4.390 ;
        RECT 15.315 1.090 15.485 4.220 ;
        RECT 15.235 0.920 15.565 1.090 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 9.835 0.920 10.165 1.090 ;
        RECT 11.995 0.920 12.325 1.090 ;
        RECT 16.315 0.920 16.645 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 9.915 0.085 10.085 0.920 ;
        RECT 12.075 0.085 12.245 0.920 ;
        RECT 16.395 0.085 16.565 0.920 ;
        RECT 0.000 -0.085 17.280 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
        RECT 10.895 -0.085 11.065 0.085 ;
        RECT 11.255 -0.085 11.425 0.085 ;
        RECT 11.615 -0.085 11.785 0.085 ;
        RECT 11.975 -0.085 12.145 0.085 ;
        RECT 12.335 -0.085 12.505 0.085 ;
        RECT 12.695 -0.085 12.865 0.085 ;
        RECT 13.055 -0.085 13.225 0.085 ;
        RECT 13.415 -0.085 13.585 0.085 ;
        RECT 13.775 -0.085 13.945 0.085 ;
        RECT 14.135 -0.085 14.305 0.085 ;
        RECT 14.495 -0.085 14.665 0.085 ;
        RECT 14.855 -0.085 15.025 0.085 ;
        RECT 15.215 -0.085 15.385 0.085 ;
        RECT 15.575 -0.085 15.745 0.085 ;
        RECT 15.935 -0.085 16.105 0.085 ;
        RECT 16.295 -0.085 16.465 0.085 ;
        RECT 16.655 -0.085 16.825 0.085 ;
        RECT 17.015 -0.085 17.185 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 17.280 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 17.280 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 9.915 5.200 10.085 6.035 ;
        RECT 12.075 5.200 12.245 6.035 ;
        RECT 16.395 5.200 16.565 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 9.835 5.030 10.165 5.200 ;
        RECT 11.995 5.030 12.325 5.200 ;
        RECT 16.315 5.030 16.645 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
        RECT 10.895 6.035 11.065 6.205 ;
        RECT 11.255 6.035 11.425 6.205 ;
        RECT 11.615 6.035 11.785 6.205 ;
        RECT 11.975 6.035 12.145 6.205 ;
        RECT 12.335 6.035 12.505 6.205 ;
        RECT 12.695 6.035 12.865 6.205 ;
        RECT 13.055 6.035 13.225 6.205 ;
        RECT 13.415 6.035 13.585 6.205 ;
        RECT 13.775 6.035 13.945 6.205 ;
        RECT 14.135 6.035 14.305 6.205 ;
        RECT 14.495 6.035 14.665 6.205 ;
        RECT 14.855 6.035 15.025 6.205 ;
        RECT 15.215 6.035 15.385 6.205 ;
        RECT 15.575 6.035 15.745 6.205 ;
        RECT 15.935 6.035 16.105 6.205 ;
        RECT 16.295 6.035 16.465 6.205 ;
        RECT 16.655 6.035 16.825 6.205 ;
        RECT 17.015 6.035 17.185 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 17.280 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 17.460 6.445 ;
      LAYER pwell ;
        RECT 0.005 1.410 1.635 1.690 ;
        RECT 5.405 1.410 7.035 1.690 ;
        RECT 9.725 1.445 11.355 1.690 ;
        RECT 8.645 1.410 11.355 1.445 ;
        RECT 15.125 1.410 16.755 1.690 ;
        RECT 0.005 0.730 16.755 1.410 ;
      LAYER li1 ;
        RECT 0.115 5.680 0.445 5.850 ;
        RECT 9.295 5.680 9.625 5.850 ;
        RECT 10.375 5.680 10.705 5.850 ;
        RECT 12.535 5.680 12.865 5.850 ;
        RECT 0.195 5.200 0.365 5.680 ;
        RECT 9.375 5.200 9.545 5.680 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 6.675 5.030 9.545 5.200 ;
        RECT 6.675 4.860 6.845 5.030 ;
        RECT 3.355 4.690 6.845 4.860 ;
        RECT 7.135 4.690 8.005 4.860 ;
        RECT 8.755 4.690 9.085 4.860 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 0.195 1.090 0.365 4.220 ;
        RECT 1.735 2.520 3.685 2.690 ;
        RECT 3.975 1.090 4.145 4.690 ;
        RECT 4.975 4.220 5.305 4.390 ;
        RECT 5.595 4.220 6.925 4.390 ;
        RECT 5.055 2.150 5.225 4.220 ;
        RECT 5.595 2.690 5.765 4.220 ;
        RECT 5.515 2.520 5.845 2.690 ;
        RECT 5.595 2.150 5.765 2.520 ;
        RECT 4.975 1.980 5.305 2.150 ;
        RECT 5.595 1.980 8.005 2.150 ;
        RECT 6.675 1.090 6.845 1.980 ;
        RECT 8.835 1.090 9.005 4.690 ;
        RECT 9.375 2.150 9.545 5.030 ;
        RECT 10.455 2.150 10.625 5.680 ;
        RECT 12.615 4.860 12.785 5.680 ;
        RECT 14.155 5.030 14.485 5.200 ;
        RECT 10.915 4.690 12.785 4.860 ;
        RECT 11.995 2.520 13.945 2.690 ;
        RECT 14.235 2.150 14.405 5.030 ;
        RECT 9.295 1.980 9.625 2.150 ;
        RECT 10.375 1.980 14.405 2.150 ;
        RECT 14.235 1.090 14.405 1.980 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 3.355 0.920 4.145 1.090 ;
        RECT 6.595 0.920 6.925 1.090 ;
        RECT 7.135 0.920 8.005 1.090 ;
        RECT 8.755 0.920 9.085 1.090 ;
        RECT 10.915 0.920 11.245 1.090 ;
        RECT 14.155 0.920 14.485 1.090 ;
        RECT 0.195 0.440 0.365 0.920 ;
        RECT 8.835 0.440 9.005 0.920 ;
        RECT 10.995 0.440 11.165 0.920 ;
        RECT 0.115 0.270 0.445 0.440 ;
        RECT 6.595 0.270 9.005 0.440 ;
        RECT 10.915 0.270 11.245 0.440 ;
  END
END DFQD1

#--------EOF---------

MACRO DFQD1_1
  CLASS CORE ;
  FOREIGN DFQD1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.200 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.166500 ;
    PORT
      LAYER li1 ;
        RECT 2.815 5.680 3.145 5.850 ;
        RECT 2.895 2.150 3.065 5.680 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END d
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.980 0.985 2.150 ;
        RECT 0.735 1.330 0.905 1.980 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 14.155 4.220 14.485 4.390 ;
        RECT 14.235 1.090 14.405 4.220 ;
        RECT 14.155 0.920 14.485 1.090 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 7.675 0.920 8.005 1.090 ;
        RECT 11.995 0.920 12.325 1.090 ;
        RECT 15.235 0.920 15.565 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 7.755 0.085 7.925 0.920 ;
        RECT 12.075 0.085 12.245 0.920 ;
        RECT 15.315 0.085 15.485 0.920 ;
        RECT 0.000 -0.085 16.200 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
        RECT 10.895 -0.085 11.065 0.085 ;
        RECT 11.255 -0.085 11.425 0.085 ;
        RECT 11.615 -0.085 11.785 0.085 ;
        RECT 11.975 -0.085 12.145 0.085 ;
        RECT 12.335 -0.085 12.505 0.085 ;
        RECT 12.695 -0.085 12.865 0.085 ;
        RECT 13.055 -0.085 13.225 0.085 ;
        RECT 13.415 -0.085 13.585 0.085 ;
        RECT 13.775 -0.085 13.945 0.085 ;
        RECT 14.135 -0.085 14.305 0.085 ;
        RECT 14.495 -0.085 14.665 0.085 ;
        RECT 14.855 -0.085 15.025 0.085 ;
        RECT 15.215 -0.085 15.385 0.085 ;
        RECT 15.575 -0.085 15.745 0.085 ;
        RECT 15.935 -0.085 16.105 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 16.200 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 16.200 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 7.755 5.200 7.925 6.035 ;
        RECT 12.075 5.200 12.245 6.035 ;
        RECT 15.315 5.200 15.485 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
        RECT 11.995 5.030 12.325 5.200 ;
        RECT 15.235 5.030 15.565 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
        RECT 10.895 6.035 11.065 6.205 ;
        RECT 11.255 6.035 11.425 6.205 ;
        RECT 11.615 6.035 11.785 6.205 ;
        RECT 11.975 6.035 12.145 6.205 ;
        RECT 12.335 6.035 12.505 6.205 ;
        RECT 12.695 6.035 12.865 6.205 ;
        RECT 13.055 6.035 13.225 6.205 ;
        RECT 13.415 6.035 13.585 6.205 ;
        RECT 13.775 6.035 13.945 6.205 ;
        RECT 14.135 6.035 14.305 6.205 ;
        RECT 14.495 6.035 14.665 6.205 ;
        RECT 14.855 6.035 15.025 6.205 ;
        RECT 15.215 6.035 15.385 6.205 ;
        RECT 15.575 6.035 15.745 6.205 ;
        RECT 15.935 6.035 16.105 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 16.200 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 16.380 6.445 ;
      LAYER pwell ;
        RECT 0.005 1.410 1.635 1.690 ;
        RECT 5.405 1.445 7.035 1.690 ;
        RECT 5.405 1.410 9.195 1.445 ;
        RECT 11.885 1.410 15.675 1.690 ;
        RECT 0.005 0.730 15.675 1.410 ;
      LAYER li1 ;
        RECT 3.355 4.690 3.685 4.860 ;
        RECT 8.295 4.690 9.085 4.860 ;
        RECT 9.835 4.690 10.165 4.860 ;
        RECT 0.115 4.220 0.905 4.390 ;
        RECT 0.735 2.690 0.905 4.220 ;
        RECT 0.195 2.520 0.985 2.690 ;
        RECT 0.195 1.090 0.365 2.520 ;
        RECT 3.435 2.150 3.605 4.690 ;
        RECT 3.895 4.220 4.225 4.390 ;
        RECT 4.435 4.220 7.465 4.390 ;
        RECT 3.975 2.690 4.145 4.220 ;
        RECT 8.295 3.230 8.465 4.690 ;
        RECT 9.915 4.390 10.085 4.690 ;
        RECT 9.915 4.220 11.165 4.390 ;
        RECT 13.075 4.220 13.405 4.390 ;
        RECT 4.975 3.060 8.465 3.230 ;
        RECT 9.295 3.060 10.625 3.230 ;
        RECT 9.375 2.690 9.545 3.060 ;
        RECT 10.455 2.690 10.625 3.060 ;
        RECT 3.895 2.520 9.545 2.690 ;
        RECT 10.375 2.520 10.705 2.690 ;
        RECT 3.435 1.980 8.545 2.150 ;
        RECT 3.435 1.090 3.605 1.980 ;
        RECT 10.995 1.500 11.165 4.220 ;
        RECT 12.535 3.060 12.865 3.230 ;
        RECT 12.615 2.150 12.785 3.060 ;
        RECT 12.535 1.980 12.865 2.150 ;
        RECT 12.615 1.500 12.785 1.980 ;
        RECT 6.675 1.330 9.545 1.500 ;
        RECT 6.675 1.090 6.845 1.330 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 6.595 0.920 6.925 1.090 ;
        RECT 8.755 0.920 9.085 1.090 ;
        RECT 8.835 0.440 9.005 0.920 ;
        RECT 9.375 0.440 9.545 1.330 ;
        RECT 9.915 1.330 12.785 1.500 ;
        RECT 9.915 1.090 10.085 1.330 ;
        RECT 13.155 1.090 13.325 4.220 ;
        RECT 9.835 0.920 10.165 1.090 ;
        RECT 13.075 0.920 13.405 1.090 ;
        RECT 13.155 0.440 13.325 0.920 ;
        RECT 8.755 0.270 9.085 0.440 ;
        RECT 9.295 0.270 9.625 0.440 ;
        RECT 13.075 0.270 13.405 0.440 ;
  END
END DFQD1_1

#--------EOF---------

MACRO DFQD1_2
  CLASS CORE ;
  FOREIGN DFQD1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.200 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.166500 ;
    PORT
      LAYER li1 ;
        RECT 4.975 3.060 5.305 3.230 ;
        RECT 5.055 2.150 5.225 3.060 ;
        RECT 4.975 1.980 5.305 2.150 ;
    END
  END d
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 14.155 4.220 14.485 4.390 ;
        RECT 14.235 1.090 14.405 4.220 ;
        RECT 14.155 0.920 14.485 1.090 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 7.675 0.920 8.005 1.090 ;
        RECT 11.995 0.920 12.325 1.090 ;
        RECT 15.235 0.920 15.565 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 7.755 0.085 7.925 0.920 ;
        RECT 12.075 0.085 12.245 0.920 ;
        RECT 15.315 0.085 15.485 0.920 ;
        RECT 0.000 -0.085 16.200 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
        RECT 10.895 -0.085 11.065 0.085 ;
        RECT 11.255 -0.085 11.425 0.085 ;
        RECT 11.615 -0.085 11.785 0.085 ;
        RECT 11.975 -0.085 12.145 0.085 ;
        RECT 12.335 -0.085 12.505 0.085 ;
        RECT 12.695 -0.085 12.865 0.085 ;
        RECT 13.055 -0.085 13.225 0.085 ;
        RECT 13.415 -0.085 13.585 0.085 ;
        RECT 13.775 -0.085 13.945 0.085 ;
        RECT 14.135 -0.085 14.305 0.085 ;
        RECT 14.495 -0.085 14.665 0.085 ;
        RECT 14.855 -0.085 15.025 0.085 ;
        RECT 15.215 -0.085 15.385 0.085 ;
        RECT 15.575 -0.085 15.745 0.085 ;
        RECT 15.935 -0.085 16.105 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 16.200 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 16.200 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 7.755 5.200 7.925 6.035 ;
        RECT 12.075 5.200 12.245 6.035 ;
        RECT 15.315 5.200 15.485 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
        RECT 11.995 5.030 12.325 5.200 ;
        RECT 15.235 5.030 15.565 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
        RECT 10.895 6.035 11.065 6.205 ;
        RECT 11.255 6.035 11.425 6.205 ;
        RECT 11.615 6.035 11.785 6.205 ;
        RECT 11.975 6.035 12.145 6.205 ;
        RECT 12.335 6.035 12.505 6.205 ;
        RECT 12.695 6.035 12.865 6.205 ;
        RECT 13.055 6.035 13.225 6.205 ;
        RECT 13.415 6.035 13.585 6.205 ;
        RECT 13.775 6.035 13.945 6.205 ;
        RECT 14.135 6.035 14.305 6.205 ;
        RECT 14.495 6.035 14.665 6.205 ;
        RECT 14.855 6.035 15.025 6.205 ;
        RECT 15.215 6.035 15.385 6.205 ;
        RECT 15.575 6.035 15.745 6.205 ;
        RECT 15.935 6.035 16.105 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 16.200 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 16.380 6.445 ;
      LAYER pwell ;
        RECT 0.005 1.410 2.715 1.690 ;
        RECT 7.565 1.410 9.195 1.445 ;
        RECT 11.885 1.410 15.675 1.690 ;
        RECT 0.005 0.730 15.675 1.410 ;
      LAYER li1 ;
        RECT 5.515 4.690 5.845 4.860 ;
        RECT 7.215 4.690 9.085 4.860 ;
        RECT 9.835 4.690 10.165 4.860 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 2.275 4.220 2.605 4.390 ;
        RECT 0.195 3.230 0.365 4.220 ;
        RECT 2.355 3.230 2.525 4.220 ;
        RECT 0.195 3.060 1.525 3.230 ;
        RECT 2.355 3.060 4.225 3.230 ;
        RECT 0.195 1.090 0.365 3.060 ;
        RECT 2.355 1.090 2.525 3.060 ;
        RECT 3.435 2.690 3.605 3.060 ;
        RECT 3.355 2.520 3.685 2.690 ;
        RECT 5.595 2.150 5.765 4.690 ;
        RECT 7.215 4.390 7.385 4.690 ;
        RECT 9.915 4.390 10.085 4.690 ;
        RECT 7.135 4.220 7.465 4.390 ;
        RECT 9.915 4.220 11.165 4.390 ;
        RECT 11.455 4.220 13.405 4.390 ;
        RECT 10.995 3.230 11.165 4.220 ;
        RECT 13.155 3.230 13.325 4.220 ;
        RECT 6.055 3.060 10.705 3.230 ;
        RECT 10.915 3.060 11.245 3.230 ;
        RECT 13.075 3.060 13.405 3.230 ;
        RECT 9.375 2.690 9.545 3.060 ;
        RECT 7.135 2.520 7.465 2.690 ;
        RECT 9.295 2.520 9.625 2.690 ;
        RECT 5.595 1.980 6.925 2.150 ;
        RECT 5.595 1.090 5.765 1.980 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 7.215 0.440 7.385 2.520 ;
        RECT 10.995 2.150 11.165 3.060 ;
        RECT 10.915 1.980 11.245 2.150 ;
        RECT 10.995 1.090 11.165 1.980 ;
        RECT 8.755 0.920 9.085 1.090 ;
        RECT 9.835 0.920 11.165 1.090 ;
        RECT 13.075 0.920 13.405 1.090 ;
        RECT 8.835 0.440 9.005 0.920 ;
        RECT 13.155 0.440 13.325 0.920 ;
        RECT 7.135 0.270 7.465 0.440 ;
        RECT 8.755 0.270 9.085 0.440 ;
        RECT 13.075 0.270 13.405 0.440 ;
  END
END DFQD1_2

#--------EOF---------

MACRO DFQD1_3
  CLASS CORE ;
  FOREIGN DFQD1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.200 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.166500 ;
    PORT
      LAYER li1 ;
        RECT 5.055 2.150 5.225 2.690 ;
        RECT 4.975 1.980 5.305 2.150 ;
    END
  END d
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.735 1.980 2.065 2.150 ;
        RECT 1.815 1.330 1.985 1.980 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 14.155 4.220 14.485 4.390 ;
        RECT 14.235 1.090 14.405 4.220 ;
        RECT 14.155 0.920 14.485 1.090 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 7.675 0.920 8.005 1.090 ;
        RECT 11.995 0.920 12.325 1.090 ;
        RECT 15.235 0.920 15.565 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 7.755 0.085 7.925 0.920 ;
        RECT 12.075 0.085 12.245 0.920 ;
        RECT 15.315 0.085 15.485 0.920 ;
        RECT 0.000 -0.085 16.200 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
        RECT 10.895 -0.085 11.065 0.085 ;
        RECT 11.255 -0.085 11.425 0.085 ;
        RECT 11.615 -0.085 11.785 0.085 ;
        RECT 11.975 -0.085 12.145 0.085 ;
        RECT 12.335 -0.085 12.505 0.085 ;
        RECT 12.695 -0.085 12.865 0.085 ;
        RECT 13.055 -0.085 13.225 0.085 ;
        RECT 13.415 -0.085 13.585 0.085 ;
        RECT 13.775 -0.085 13.945 0.085 ;
        RECT 14.135 -0.085 14.305 0.085 ;
        RECT 14.495 -0.085 14.665 0.085 ;
        RECT 14.855 -0.085 15.025 0.085 ;
        RECT 15.215 -0.085 15.385 0.085 ;
        RECT 15.575 -0.085 15.745 0.085 ;
        RECT 15.935 -0.085 16.105 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 16.200 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 16.200 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 7.755 5.200 7.925 6.035 ;
        RECT 12.075 5.200 12.245 6.035 ;
        RECT 15.315 5.200 15.485 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
        RECT 11.995 5.030 12.325 5.200 ;
        RECT 15.235 5.030 15.565 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
        RECT 10.895 6.035 11.065 6.205 ;
        RECT 11.255 6.035 11.425 6.205 ;
        RECT 11.615 6.035 11.785 6.205 ;
        RECT 11.975 6.035 12.145 6.205 ;
        RECT 12.335 6.035 12.505 6.205 ;
        RECT 12.695 6.035 12.865 6.205 ;
        RECT 13.055 6.035 13.225 6.205 ;
        RECT 13.415 6.035 13.585 6.205 ;
        RECT 13.775 6.035 13.945 6.205 ;
        RECT 14.135 6.035 14.305 6.205 ;
        RECT 14.495 6.035 14.665 6.205 ;
        RECT 14.855 6.035 15.025 6.205 ;
        RECT 15.215 6.035 15.385 6.205 ;
        RECT 15.575 6.035 15.745 6.205 ;
        RECT 15.935 6.035 16.105 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 16.200 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 16.380 6.445 ;
      LAYER pwell ;
        RECT 0.005 1.410 2.715 1.690 ;
        RECT 7.565 1.410 9.195 1.445 ;
        RECT 11.885 1.410 15.675 1.690 ;
        RECT 0.005 0.730 15.675 1.410 ;
      LAYER li1 ;
        RECT 9.375 5.680 10.705 5.850 ;
        RECT 5.515 4.690 5.845 4.860 ;
        RECT 8.755 4.690 9.085 4.860 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 2.275 4.220 3.145 4.390 ;
        RECT 0.195 3.230 0.365 4.220 ;
        RECT 5.595 3.230 5.765 4.690 ;
        RECT 0.195 3.060 4.225 3.230 ;
        RECT 5.595 3.060 8.005 3.230 ;
        RECT 0.195 1.090 0.365 3.060 ;
        RECT 1.195 2.520 4.225 2.690 ;
        RECT 2.355 1.090 2.525 2.520 ;
        RECT 5.595 1.090 5.765 3.060 ;
        RECT 8.835 2.150 9.005 4.690 ;
        RECT 9.375 2.150 9.545 5.680 ;
        RECT 9.835 4.690 10.165 4.860 ;
        RECT 9.915 3.230 10.085 4.690 ;
        RECT 13.075 4.220 13.405 4.390 ;
        RECT 9.915 3.060 12.865 3.230 ;
        RECT 7.135 1.980 9.005 2.150 ;
        RECT 9.295 1.980 9.625 2.150 ;
        RECT 8.835 1.090 9.005 1.980 ;
        RECT 9.915 1.090 10.085 3.060 ;
        RECT 12.615 2.150 12.785 3.060 ;
        RECT 12.535 1.980 12.865 2.150 ;
        RECT 13.155 1.090 13.325 4.220 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 8.755 0.920 9.085 1.090 ;
        RECT 9.835 0.920 10.165 1.090 ;
        RECT 13.075 0.920 13.405 1.090 ;
        RECT 0.195 0.440 0.365 0.920 ;
        RECT 13.155 0.440 13.325 0.920 ;
        RECT 0.115 0.270 0.445 0.440 ;
        RECT 13.075 0.270 13.405 0.440 ;
  END
END DFQD1_3

#--------EOF---------

MACRO FILL1
  CLASS CORE ;
  FOREIGN FILL1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.360 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 0.360 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 0.360 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 0.360 6.205 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 0.360 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 0.540 6.445 ;
  END
END FILL1

#--------EOF---------

MACRO FILL2
  CLASS CORE ;
  FOREIGN FILL2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.720 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 0.720 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 0.720 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 0.720 6.205 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 0.720 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 0.900 6.445 ;
  END
END FILL2

#--------EOF---------

MACRO FILL4
  CLASS CORE ;
  FOREIGN FILL4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.440 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 1.440 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 1.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 1.440 6.205 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 1.440 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 1.620 6.445 ;
  END
END FILL4

#--------EOF---------

MACRO FILL8
  CLASS CORE ;
  FOREIGN FILL8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.880 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 2.880 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 2.880 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 2.880 6.205 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 2.880 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 3.060 6.445 ;
  END
END FILL8

#--------EOF---------

MACRO INVD1
  CLASS CORE ;
  FOREIGN INVD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.160 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 0.195 1.090 0.365 4.220 ;
        RECT 0.115 0.920 0.445 1.090 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 0.000 -0.085 2.160 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 2.160 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 2.160 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 2.160 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 2.340 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 1.635 1.690 ;
  END
END INVD1

#--------EOF---------

MACRO MUX2D1
  CLASS CORE ;
  FOREIGN MUX2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.291000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 0.440 0.905 1.090 ;
        RECT 0.655 0.270 0.985 0.440 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.735 1.980 2.065 2.150 ;
        RECT 1.815 1.330 1.985 1.980 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.212250 ;
    PORT
      LAYER li1 ;
        RECT 2.815 1.980 3.145 2.150 ;
        RECT 2.895 1.330 3.065 1.980 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.896700 ;
    PORT
      LAYER li1 ;
        RECT 7.675 4.690 8.005 4.860 ;
        RECT 7.755 1.090 7.925 4.690 ;
        RECT 7.675 0.920 8.005 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 6.595 0.920 6.925 1.090 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 6.675 0.085 6.845 0.920 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.640 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 8.640 6.205 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 6.675 5.200 6.845 6.035 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 6.595 5.030 6.925 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 8.640 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 8.820 6.445 ;
      LAYER pwell ;
        RECT 1.085 1.495 2.715 1.690 ;
        RECT 1.085 1.410 3.795 1.495 ;
        RECT 6.485 1.410 8.115 1.690 ;
        RECT 0.005 0.730 8.115 1.410 ;
      LAYER li1 ;
        RECT 3.355 5.680 5.765 5.850 ;
        RECT 5.595 5.200 5.765 5.680 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 4.435 5.030 5.305 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 0.195 2.690 0.365 5.030 ;
        RECT 3.355 4.690 3.685 4.860 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 1.275 3.230 1.445 4.220 ;
        RECT 3.435 3.230 3.605 4.690 ;
        RECT 1.195 3.060 1.525 3.230 ;
        RECT 3.355 3.060 3.685 3.230 ;
        RECT 4.515 2.690 4.685 5.030 ;
        RECT 5.595 3.230 5.765 5.030 ;
        RECT 5.515 3.060 5.845 3.230 ;
        RECT 0.195 2.520 4.685 2.690 ;
        RECT 0.195 1.090 0.365 2.520 ;
        RECT 1.195 1.980 1.525 2.150 ;
        RECT 3.355 1.980 3.685 2.150 ;
        RECT 1.275 1.090 1.445 1.980 ;
        RECT 3.435 1.090 3.605 1.980 ;
        RECT 4.515 1.090 4.685 2.520 ;
        RECT 5.595 1.090 5.765 3.060 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
  END
END MUX2D1

#--------EOF---------

MACRO MUX2D1_1
  CLASS CORE ;
  FOREIGN MUX2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.291000 ;
    PORT
      LAYER li1 ;
        RECT 1.735 5.680 2.065 5.850 ;
        RECT 1.815 2.690 1.985 5.680 ;
        RECT 1.735 2.520 2.065 2.690 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.212250 ;
    PORT
      LAYER li1 ;
        RECT 3.895 2.520 4.685 2.690 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.896700 ;
    PORT
      LAYER li1 ;
        RECT 6.595 4.690 6.925 4.860 ;
        RECT 6.675 1.090 6.845 4.690 ;
        RECT 6.595 0.920 6.925 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 7.675 0.920 8.005 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 7.755 0.085 7.925 0.920 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.640 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 8.640 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 7.755 5.200 7.925 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 8.640 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 8.820 6.445 ;
      LAYER pwell ;
        RECT 0.005 1.410 1.635 1.690 ;
        RECT 3.245 1.410 4.875 1.495 ;
        RECT 6.485 1.410 8.115 1.690 ;
        RECT 0.005 0.730 8.115 1.410 ;
      LAYER li1 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 5.055 5.030 5.845 5.200 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 1.275 1.090 1.445 4.220 ;
        RECT 2.355 1.090 2.525 5.030 ;
        RECT 2.895 4.690 3.685 4.860 ;
        RECT 2.895 1.090 3.065 4.690 ;
        RECT 5.055 3.230 5.225 5.030 ;
        RECT 3.355 3.060 5.225 3.230 ;
        RECT 3.355 1.980 5.765 2.150 ;
        RECT 5.595 1.090 5.765 1.980 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 2.895 0.920 3.685 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 2.355 0.440 2.525 0.920 ;
        RECT 2.275 0.270 2.605 0.440 ;
  END
END MUX2D1_1

#--------EOF---------

MACRO MUX2D1_2
  CLASS CORE ;
  FOREIGN MUX2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.291000 ;
    PORT
      LAYER li1 ;
        RECT 3.895 1.980 4.685 2.150 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.815 1.980 3.145 2.150 ;
        RECT 2.895 1.330 3.065 1.980 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.212250 ;
    PORT
      LAYER li1 ;
        RECT 1.735 1.980 2.065 2.150 ;
        RECT 1.815 1.330 1.985 1.980 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.896700 ;
    PORT
      LAYER li1 ;
        RECT 7.675 4.690 8.005 4.860 ;
        RECT 7.755 1.090 7.925 4.690 ;
        RECT 7.675 0.920 8.005 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 6.595 0.920 6.925 1.090 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 6.675 0.085 6.845 0.920 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.640 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 8.640 6.205 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 6.675 5.200 6.845 6.035 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 6.595 5.030 6.925 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 8.640 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 8.820 6.445 ;
      LAYER pwell ;
        RECT 2.165 1.495 3.795 1.690 ;
        RECT 1.085 1.410 3.795 1.495 ;
        RECT 6.485 1.410 8.115 1.690 ;
        RECT 0.005 0.730 8.115 1.410 ;
      LAYER li1 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
        RECT 5.055 5.030 5.845 5.200 ;
        RECT 0.195 2.690 0.365 5.030 ;
        RECT 1.195 4.690 1.525 4.860 ;
        RECT 1.275 3.230 1.445 4.690 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 3.435 3.230 3.605 4.220 ;
        RECT 1.195 3.060 1.525 3.230 ;
        RECT 3.355 3.060 3.685 3.230 ;
        RECT 4.515 2.690 4.685 5.030 ;
        RECT 5.055 4.390 5.225 5.030 ;
        RECT 4.975 4.220 5.305 4.390 ;
        RECT 0.195 2.520 4.765 2.690 ;
        RECT 0.195 1.090 0.365 2.520 ;
        RECT 1.195 1.980 1.525 2.150 ;
        RECT 3.355 1.980 3.685 2.150 ;
        RECT 1.275 1.090 1.445 1.980 ;
        RECT 3.435 1.090 3.605 1.980 ;
        RECT 5.055 1.500 5.225 4.220 ;
        RECT 3.975 1.330 5.765 1.500 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 3.975 0.440 4.145 1.330 ;
        RECT 5.595 1.090 5.765 1.330 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 4.515 0.440 4.685 0.920 ;
        RECT 3.895 0.270 4.225 0.440 ;
        RECT 4.435 0.270 4.765 0.440 ;
  END
END MUX2D1_2

#--------EOF---------

MACRO MUX2D1_3
  CLASS CORE ;
  FOREIGN MUX2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.291000 ;
    PORT
      LAYER li1 ;
        RECT 1.735 5.680 3.065 5.850 ;
        RECT 2.895 4.860 3.065 5.680 ;
        RECT 2.895 4.690 5.225 4.860 ;
        RECT 2.895 3.230 3.065 4.690 ;
        RECT 5.055 4.390 5.225 4.690 ;
        RECT 4.975 4.220 5.305 4.390 ;
        RECT 2.815 3.060 3.145 3.230 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 3.895 1.980 4.225 2.150 ;
        RECT 3.975 1.330 4.145 1.980 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.212250 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.896700 ;
    PORT
      LAYER li1 ;
        RECT 6.595 4.690 6.925 4.860 ;
        RECT 6.675 1.090 6.845 4.690 ;
        RECT 6.595 0.920 6.925 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 7.675 0.920 8.005 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 7.755 0.085 7.925 0.920 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.640 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 8.640 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 7.755 5.200 7.925 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 8.640 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 8.820 6.445 ;
      LAYER pwell ;
        RECT 0.005 1.410 1.635 1.495 ;
        RECT 3.245 1.410 4.875 1.690 ;
        RECT 6.485 1.410 8.115 1.690 ;
        RECT 0.005 0.730 8.115 1.410 ;
      LAYER li1 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 5.515 5.030 6.305 5.200 ;
        RECT 1.195 4.690 1.525 4.860 ;
        RECT 1.275 1.090 1.445 4.690 ;
        RECT 2.355 2.690 2.525 5.030 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 3.435 3.230 3.605 4.220 ;
        RECT 3.355 3.060 3.685 3.230 ;
        RECT 2.355 2.520 5.845 2.690 ;
        RECT 2.355 1.090 2.525 2.520 ;
        RECT 3.355 1.980 3.685 2.150 ;
        RECT 3.435 1.090 3.605 1.980 ;
        RECT 6.135 1.090 6.305 5.030 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 5.515 0.920 6.305 1.090 ;
        RECT 5.595 0.440 5.765 0.920 ;
        RECT 5.515 0.270 5.845 0.440 ;
  END
END MUX2D1_3

#--------EOF---------

MACRO ND2D1
  CLASS CORE ;
  FOREIGN ND2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.450000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 1.275 3.230 1.445 4.220 ;
        RECT 1.275 3.060 2.525 3.230 ;
        RECT 2.355 1.090 2.525 3.060 ;
        RECT 2.275 0.920 2.605 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 0.000 -0.085 3.240 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.240 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 3.240 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 3.240 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 3.420 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 2.715 1.690 ;
  END
END ND2D1

#--------EOF---------

MACRO ND2D1_1
  CLASS CORE ;
  FOREIGN ND2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.450000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 1.275 3.230 1.445 4.220 ;
        RECT 0.195 3.060 1.445 3.230 ;
        RECT 0.195 1.090 0.365 3.060 ;
        RECT 0.115 0.920 0.445 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 0.000 -0.085 3.240 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.240 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 3.240 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 3.240 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 3.420 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 2.715 1.690 ;
  END
END ND2D1_1

#--------EOF---------

MACRO ND2D1_2
  CLASS CORE ;
  FOREIGN ND2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.769000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 4.690 2.605 4.860 ;
        RECT 2.275 4.220 2.605 4.390 ;
        RECT 2.355 1.090 2.525 4.220 ;
        RECT 2.275 0.920 2.605 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 0.000 -0.085 3.240 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.240 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 3.240 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 3.240 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 3.420 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 2.715 1.690 ;
  END
END ND2D1_2

#--------EOF---------

MACRO ND2D1_3
  CLASS CORE ;
  FOREIGN ND2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.769000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 4.690 2.605 4.860 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 0.195 1.090 0.365 4.220 ;
        RECT 0.115 0.920 0.445 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 0.000 -0.085 3.240 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.240 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 3.240 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 3.240 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 3.420 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 2.715 1.690 ;
  END
END ND2D1_3

#--------EOF---------

MACRO ND3D1
  CLASS CORE ;
  FOREIGN ND3D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.121000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 1.275 3.230 1.445 4.220 ;
        RECT 3.435 3.230 3.605 4.220 ;
        RECT 0.195 3.060 3.605 3.230 ;
        RECT 0.195 1.090 0.365 3.060 ;
        RECT 0.115 0.920 0.445 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.320 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 4.320 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 4.320 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 4.500 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 3.795 1.690 ;
  END
END ND3D1

#--------EOF---------

MACRO ND3D1_1
  CLASS CORE ;
  FOREIGN ND3D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.121000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 1.275 1.090 1.445 4.220 ;
        RECT 3.435 1.500 3.605 4.220 ;
        RECT 2.355 1.330 3.605 1.500 ;
        RECT 2.355 1.090 2.525 1.330 ;
        RECT 1.275 0.920 2.605 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 3.975 2.150 4.145 2.690 ;
        RECT 3.895 1.980 4.225 2.150 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 5.400 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.400 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 5.400 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 5.400 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 5.580 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 4.875 1.690 ;
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 0.195 0.440 0.365 0.920 ;
        RECT 3.435 0.440 3.605 0.920 ;
        RECT 0.195 0.270 3.605 0.440 ;
  END
END ND3D1_1

#--------EOF---------

MACRO ND3D1_2
  CLASS CORE ;
  FOREIGN ND3D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.121000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 1.275 2.150 1.445 4.220 ;
        RECT 3.435 2.150 3.605 4.220 ;
        RECT 1.275 1.980 3.605 2.150 ;
        RECT 3.435 1.090 3.605 1.980 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.690 3.065 3.230 ;
        RECT 2.815 2.520 3.145 2.690 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.690 1.985 3.230 ;
        RECT 1.735 2.520 2.065 2.690 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.320 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 4.320 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 4.320 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 4.500 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 3.795 1.690 ;
  END
END ND3D1_2

#--------EOF---------

MACRO ND3D1_3
  CLASS CORE ;
  FOREIGN ND3D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.121000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 5.030 1.525 5.200 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 1.275 3.230 1.445 4.220 ;
        RECT 1.275 3.060 2.525 3.230 ;
        RECT 2.355 2.150 2.525 3.060 ;
        RECT 3.435 2.150 3.605 4.220 ;
        RECT 2.355 1.980 3.605 2.150 ;
        RECT 3.435 1.090 3.605 1.980 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 3.975 2.150 4.145 2.690 ;
        RECT 3.895 1.980 4.225 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 0.000 -0.085 5.400 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.400 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 5.400 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 5.400 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 5.580 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 4.875 1.690 ;
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 3.975 0.920 4.765 1.090 ;
        RECT 0.195 0.440 0.365 0.920 ;
        RECT 3.975 0.440 4.145 0.920 ;
        RECT 0.115 0.270 0.445 0.440 ;
        RECT 2.815 0.270 4.145 0.440 ;
  END
END ND3D1_3

#--------EOF---------

MACRO ND4D1
  CLASS CORE ;
  FOREIGN ND4D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 5.055 2.150 5.225 2.690 ;
        RECT 4.975 1.980 5.305 2.150 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a3
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.792000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 4.435 4.220 4.765 4.390 ;
        RECT 1.275 3.230 1.445 4.220 ;
        RECT 3.435 3.230 3.605 4.220 ;
        RECT 4.515 3.230 4.685 4.220 ;
        RECT 1.275 3.060 4.685 3.230 ;
        RECT 3.435 1.090 3.605 3.060 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 0.000 -0.085 6.480 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.480 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 6.480 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 6.480 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 6.660 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 5.955 1.690 ;
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 0.195 0.440 0.365 0.920 ;
        RECT 4.515 0.440 4.685 0.920 ;
        RECT 0.195 0.270 4.685 0.440 ;
  END
END ND4D1

#--------EOF---------

MACRO ND4D1_1
  CLASS CORE ;
  FOREIGN ND4D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a3
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.792000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 4.765 4.390 ;
        RECT 4.515 1.090 4.685 4.220 ;
        RECT 4.435 0.920 4.765 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 5.055 2.150 5.225 2.690 ;
        RECT 4.975 1.980 5.305 2.150 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 0.000 -0.085 6.480 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.480 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 6.480 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 6.480 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 6.660 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 5.955 1.690 ;
      LAYER li1 ;
        RECT 2.895 1.330 4.145 1.500 ;
        RECT 2.895 1.090 3.065 1.330 ;
        RECT 0.115 0.920 3.065 1.090 ;
        RECT 3.975 0.440 4.145 1.330 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 5.595 0.440 5.765 0.920 ;
        RECT 3.975 0.270 5.765 0.440 ;
  END
END ND4D1_1

#--------EOF---------

MACRO ND4D1_2
  CLASS CORE ;
  FOREIGN ND4D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.815 5.680 3.145 5.850 ;
        RECT 2.895 2.690 3.065 5.680 ;
        RECT 2.815 2.520 3.145 2.690 ;
    END
  END a2
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.735 5.680 2.065 5.850 ;
        RECT 1.815 2.150 1.985 5.680 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a3
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.473000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 1.275 1.090 1.445 4.220 ;
        RECT 3.435 1.090 3.605 4.220 ;
        RECT 1.275 0.920 4.765 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 3.975 2.150 4.145 2.690 ;
        RECT 3.895 1.980 4.225 2.150 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 0.000 -0.085 5.400 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.400 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 5.400 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 5.400 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 5.580 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 4.875 1.690 ;
  END
END ND4D1_2

#--------EOF---------

MACRO ND4D1_3
  CLASS CORE ;
  FOREIGN ND4D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 3.975 2.150 4.145 2.690 ;
        RECT 3.895 1.980 4.225 2.150 ;
    END
  END a2
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.735 5.680 2.065 5.850 ;
        RECT 1.815 2.690 1.985 5.680 ;
        RECT 1.735 2.520 2.065 2.690 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a3
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.473000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 4.435 4.220 4.765 4.390 ;
        RECT 1.275 1.500 1.445 4.220 ;
        RECT 4.515 1.500 4.685 4.220 ;
        RECT 1.275 1.330 5.765 1.500 ;
        RECT 5.595 1.090 5.765 1.330 ;
        RECT 5.515 0.920 5.845 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 5.055 2.150 5.225 2.690 ;
        RECT 4.975 1.980 5.305 2.150 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 0.000 -0.085 6.480 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.480 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 6.480 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 6.480 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 6.660 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 5.955 1.690 ;
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 0.195 0.440 0.365 0.920 ;
        RECT 3.435 0.440 3.605 0.920 ;
        RECT 0.115 0.270 0.445 0.440 ;
        RECT 3.355 0.270 3.685 0.440 ;
  END
END ND4D1_3

#--------EOF---------

MACRO NR2D1
  CLASS CORE ;
  FOREIGN NR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.322000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 4.220 1.445 4.390 ;
        RECT 1.275 1.090 1.445 4.220 ;
        RECT 1.195 0.920 1.525 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 0.000 -0.085 3.240 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.240 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 3.240 6.205 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 2.275 5.030 2.605 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 3.240 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 3.420 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 2.715 1.690 ;
  END
END NR2D1

#--------EOF---------

MACRO NR2D1_1
  CLASS CORE ;
  FOREIGN NR2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.322000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 4.220 2.605 4.390 ;
        RECT 2.355 3.230 2.525 4.220 ;
        RECT 1.275 3.060 2.525 3.230 ;
        RECT 1.275 1.090 1.445 3.060 ;
        RECT 1.195 0.920 1.525 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 0.000 -0.085 3.240 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.240 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 3.240 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 3.240 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 3.420 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 2.715 1.690 ;
  END
END NR2D1_1

#--------EOF---------

MACRO NR2D1_2
  CLASS CORE ;
  FOREIGN NR2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.525000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 0.195 1.500 0.365 4.220 ;
        RECT 0.195 1.330 2.525 1.500 ;
        RECT 0.195 1.090 0.365 1.330 ;
        RECT 2.355 1.090 2.525 1.330 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 0.000 -0.085 3.240 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.240 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 3.240 6.205 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 2.275 5.030 2.605 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 3.240 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 3.420 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 2.715 1.690 ;
  END
END NR2D1_2

#--------EOF---------

MACRO NR2D1_3
  CLASS CORE ;
  FOREIGN NR2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.240 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.525000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 4.220 2.605 4.390 ;
        RECT 0.195 1.330 1.985 1.500 ;
        RECT 0.195 1.090 0.365 1.330 ;
        RECT 1.815 1.090 1.985 1.330 ;
        RECT 2.355 1.090 2.525 4.220 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 1.815 0.920 2.605 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 0.000 -0.085 3.240 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.240 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 3.240 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 3.240 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 3.420 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 2.715 1.690 ;
  END
END NR2D1_3

#--------EOF---------

MACRO NR3D1
  CLASS CORE ;
  FOREIGN NR3D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.800 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.101000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 4.220 1.525 4.390 ;
        RECT 0.735 1.090 0.905 4.220 ;
        RECT 1.275 1.330 3.605 1.500 ;
        RECT 1.275 1.090 1.445 1.330 ;
        RECT 3.435 1.090 3.605 1.330 ;
        RECT 0.735 0.920 1.525 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 4.975 3.060 5.305 3.230 ;
        RECT 5.055 2.150 5.225 3.060 ;
        RECT 1.195 1.980 5.225 2.150 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 5.595 2.150 5.765 2.690 ;
        RECT 5.515 1.980 5.845 2.150 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.690 1.985 3.230 ;
        RECT 1.735 2.520 2.065 2.690 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 0.000 -0.085 10.800 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 10.800 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 10.800 6.205 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 7.755 5.200 7.925 6.035 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 10.800 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 10.980 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 3.795 1.690 ;
      LAYER li1 ;
        RECT 0.115 4.690 9.085 4.860 ;
        RECT 3.355 4.220 4.765 4.390 ;
        RECT 6.595 4.220 10.165 4.390 ;
  END
END NR3D1

#--------EOF---------

MACRO NR3D1_1
  CLASS CORE ;
  FOREIGN NR3D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.880 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.101000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 1.275 1.500 1.445 4.220 ;
        RECT 1.275 1.330 3.605 1.500 ;
        RECT 1.275 1.090 1.445 1.330 ;
        RECT 3.435 1.090 3.605 1.330 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 6.055 3.060 6.385 3.230 ;
        RECT 6.135 2.690 6.305 3.060 ;
        RECT 1.735 2.520 6.305 2.690 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 3.895 1.980 4.225 2.150 ;
        RECT 3.975 1.330 4.145 1.980 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 0.655 5.680 0.985 5.850 ;
        RECT 0.735 2.690 0.905 5.680 ;
        RECT 0.655 2.520 0.985 2.690 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 11.880 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
        RECT 10.895 -0.085 11.065 0.085 ;
        RECT 11.255 -0.085 11.425 0.085 ;
        RECT 11.615 -0.085 11.785 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 11.880 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 11.880 6.205 ;
        RECT 6.675 5.200 6.845 6.035 ;
        RECT 8.835 5.200 9.005 6.035 ;
        RECT 6.595 5.030 6.925 5.200 ;
        RECT 8.755 5.030 9.085 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
        RECT 10.895 6.035 11.065 6.205 ;
        RECT 11.255 6.035 11.425 6.205 ;
        RECT 11.615 6.035 11.785 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 11.880 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 12.060 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 4.875 1.690 ;
      LAYER li1 ;
        RECT 2.275 4.690 10.165 4.860 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 4.435 4.220 5.845 4.390 ;
        RECT 7.675 4.220 11.245 4.390 ;
        RECT 0.195 3.230 0.365 4.220 ;
        RECT 3.435 3.230 3.605 4.220 ;
        RECT 0.115 3.060 0.445 3.230 ;
        RECT 3.355 3.060 3.685 3.230 ;
  END
END NR3D1_1

#--------EOF---------

MACRO NR3D1_2
  CLASS CORE ;
  FOREIGN NR3D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.800 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.101000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 1.275 3.230 1.445 4.220 ;
        RECT 0.195 3.060 1.445 3.230 ;
        RECT 0.195 1.500 0.365 3.060 ;
        RECT 0.195 1.330 2.525 1.500 ;
        RECT 0.195 1.090 0.365 1.330 ;
        RECT 2.355 1.090 2.525 1.330 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 0.440 0.905 1.090 ;
        RECT 0.655 0.270 0.985 0.440 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 2.815 3.060 9.625 3.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 0.000 -0.085 10.800 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 10.800 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 10.800 6.205 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 7.755 5.200 7.925 6.035 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 10.800 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 10.980 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 3.795 1.690 ;
      LAYER li1 ;
        RECT 0.115 4.690 9.085 4.860 ;
        RECT 3.355 4.220 4.765 4.390 ;
        RECT 6.595 4.220 10.165 4.390 ;
  END
END NR3D1_2

#--------EOF---------

MACRO NR3D1_3
  CLASS CORE ;
  FOREIGN NR3D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.800 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.101000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 4.220 2.605 4.390 ;
        RECT 2.355 3.230 2.525 4.220 ;
        RECT 2.355 3.060 3.605 3.230 ;
        RECT 3.435 1.500 3.605 3.060 ;
        RECT 1.275 1.330 3.605 1.500 ;
        RECT 1.275 1.090 1.445 1.330 ;
        RECT 3.435 1.090 3.605 1.330 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 0.655 5.680 0.985 5.850 ;
        RECT 0.735 2.690 0.905 5.680 ;
        RECT 0.655 2.520 0.985 2.690 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 1.735 5.680 3.145 5.850 ;
        RECT 1.815 2.690 1.985 5.680 ;
        RECT 1.735 2.520 2.065 2.690 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 0.000 -0.085 10.800 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 10.800 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 10.800 6.205 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 7.755 5.200 7.925 6.035 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 10.800 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 10.980 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 3.795 1.690 ;
      LAYER li1 ;
        RECT 3.355 4.690 9.085 4.860 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 4.435 4.220 4.765 4.390 ;
        RECT 6.595 4.220 10.165 4.390 ;
        RECT 0.195 3.230 0.365 4.220 ;
        RECT 4.515 3.230 4.685 4.220 ;
        RECT 0.115 3.060 0.445 3.230 ;
        RECT 4.435 3.060 4.765 3.230 ;
  END
END NR3D1_3

#--------EOF---------

MACRO NR4D1
  CLASS CORE ;
  FOREIGN NR4D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.869300 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 1.985 4.390 ;
        RECT 1.815 2.150 1.985 4.220 ;
        RECT 1.275 1.980 4.685 2.150 ;
        RECT 1.275 1.090 1.445 1.980 ;
        RECT 4.515 1.090 4.685 1.980 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
    END
  END zn
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 5.055 2.150 5.225 2.690 ;
        RECT 4.975 1.980 5.305 2.150 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 3.975 0.440 4.145 1.090 ;
        RECT 3.895 0.270 4.225 0.440 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.690 3.065 3.230 ;
        RECT 2.815 2.520 3.145 2.690 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 0.655 3.060 0.985 3.230 ;
        RECT 0.735 0.440 0.905 3.060 ;
        RECT 0.655 0.270 0.985 0.440 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 0.000 -0.085 15.120 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
        RECT 10.895 -0.085 11.065 0.085 ;
        RECT 11.255 -0.085 11.425 0.085 ;
        RECT 11.615 -0.085 11.785 0.085 ;
        RECT 11.975 -0.085 12.145 0.085 ;
        RECT 12.335 -0.085 12.505 0.085 ;
        RECT 12.695 -0.085 12.865 0.085 ;
        RECT 13.055 -0.085 13.225 0.085 ;
        RECT 13.415 -0.085 13.585 0.085 ;
        RECT 13.775 -0.085 13.945 0.085 ;
        RECT 14.135 -0.085 14.305 0.085 ;
        RECT 14.495 -0.085 14.665 0.085 ;
        RECT 14.855 -0.085 15.025 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 15.120 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 15.120 6.205 ;
        RECT 9.915 5.200 10.085 6.035 ;
        RECT 12.075 5.200 12.245 6.035 ;
        RECT 9.835 5.030 10.165 5.200 ;
        RECT 11.995 5.030 12.325 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
        RECT 10.895 6.035 11.065 6.205 ;
        RECT 11.255 6.035 11.425 6.205 ;
        RECT 11.615 6.035 11.785 6.205 ;
        RECT 11.975 6.035 12.145 6.205 ;
        RECT 12.335 6.035 12.505 6.205 ;
        RECT 12.695 6.035 12.865 6.205 ;
        RECT 13.055 6.035 13.225 6.205 ;
        RECT 13.415 6.035 13.585 6.205 ;
        RECT 13.775 6.035 13.945 6.205 ;
        RECT 14.135 6.035 14.305 6.205 ;
        RECT 14.495 6.035 14.665 6.205 ;
        RECT 14.855 6.035 15.025 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 15.120 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 15.300 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 5.955 1.445 ;
      LAYER li1 ;
        RECT 0.115 4.690 3.685 4.860 ;
        RECT 5.515 4.690 8.465 4.860 ;
        RECT 8.755 4.690 14.485 4.860 ;
        RECT 8.295 4.390 8.465 4.690 ;
        RECT 2.275 4.220 6.925 4.390 ;
        RECT 7.675 4.220 8.005 4.390 ;
        RECT 8.295 4.220 11.245 4.390 ;
        RECT 13.075 4.220 13.405 4.390 ;
        RECT 7.755 3.230 7.925 4.220 ;
        RECT 13.155 3.230 13.325 4.220 ;
        RECT 7.755 3.060 13.325 3.230 ;
  END
END NR4D1

#--------EOF---------

MACRO NR4D1_1
  CLASS CORE ;
  FOREIGN NR4D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.040 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.869300 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 1.275 1.500 1.445 4.220 ;
        RECT 1.275 1.330 3.605 1.500 ;
        RECT 1.275 1.090 1.445 1.330 ;
        RECT 3.435 1.090 3.605 1.330 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END zn
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 4.515 2.150 4.685 2.690 ;
        RECT 4.435 1.980 4.765 2.150 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 3.895 3.060 4.225 3.230 ;
        RECT 3.975 0.440 4.145 3.060 ;
        RECT 3.895 0.270 4.225 0.440 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 14.040 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
        RECT 10.895 -0.085 11.065 0.085 ;
        RECT 11.255 -0.085 11.425 0.085 ;
        RECT 11.615 -0.085 11.785 0.085 ;
        RECT 11.975 -0.085 12.145 0.085 ;
        RECT 12.335 -0.085 12.505 0.085 ;
        RECT 12.695 -0.085 12.865 0.085 ;
        RECT 13.055 -0.085 13.225 0.085 ;
        RECT 13.415 -0.085 13.585 0.085 ;
        RECT 13.775 -0.085 13.945 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 14.040 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 14.040 6.205 ;
        RECT 8.835 5.200 9.005 6.035 ;
        RECT 10.995 5.200 11.165 6.035 ;
        RECT 8.755 5.030 9.085 5.200 ;
        RECT 10.915 5.030 11.245 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
        RECT 10.895 6.035 11.065 6.205 ;
        RECT 11.255 6.035 11.425 6.205 ;
        RECT 11.615 6.035 11.785 6.205 ;
        RECT 11.975 6.035 12.145 6.205 ;
        RECT 12.335 6.035 12.505 6.205 ;
        RECT 12.695 6.035 12.865 6.205 ;
        RECT 13.055 6.035 13.225 6.205 ;
        RECT 13.415 6.035 13.585 6.205 ;
        RECT 13.775 6.035 13.945 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 14.040 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 14.220 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 4.875 1.445 ;
      LAYER li1 ;
        RECT 0.115 5.030 5.845 5.200 ;
        RECT 4.435 4.690 7.385 4.860 ;
        RECT 7.675 4.690 13.405 4.860 ;
        RECT 7.215 4.390 7.385 4.690 ;
        RECT 6.595 4.220 6.925 4.390 ;
        RECT 7.215 4.220 10.165 4.390 ;
        RECT 11.995 4.220 12.325 4.390 ;
        RECT 6.675 3.230 6.845 4.220 ;
        RECT 12.075 3.230 12.245 4.220 ;
        RECT 6.675 3.060 12.245 3.230 ;
  END
END NR4D1_1

#--------EOF---------

MACRO NR4D1_2
  CLASS CORE ;
  FOREIGN NR4D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.120 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.869300 ;
    PORT
      LAYER li1 ;
        RECT 3.975 4.220 4.765 4.390 ;
        RECT 3.975 1.500 4.145 4.220 ;
        RECT 1.275 1.330 4.145 1.500 ;
        RECT 1.275 1.090 1.445 1.330 ;
        RECT 3.975 1.090 4.145 1.330 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 3.975 0.920 4.765 1.090 ;
    END
  END zn
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.690 1.985 3.230 ;
        RECT 1.735 2.520 2.065 2.690 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 0.735 0.440 0.905 1.090 ;
        RECT 0.655 0.270 0.985 0.440 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 0.655 3.060 0.985 3.230 ;
        RECT 7.135 3.060 7.465 3.230 ;
        RECT 0.735 2.150 0.905 3.060 ;
        RECT 7.215 2.150 7.385 3.060 ;
        RECT 0.735 1.980 3.145 2.150 ;
        RECT 4.435 1.980 7.385 2.150 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 5.055 2.690 5.225 3.230 ;
        RECT 4.975 2.520 5.305 2.690 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 0.000 -0.085 15.120 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
        RECT 10.895 -0.085 11.065 0.085 ;
        RECT 11.255 -0.085 11.425 0.085 ;
        RECT 11.615 -0.085 11.785 0.085 ;
        RECT 11.975 -0.085 12.145 0.085 ;
        RECT 12.335 -0.085 12.505 0.085 ;
        RECT 12.695 -0.085 12.865 0.085 ;
        RECT 13.055 -0.085 13.225 0.085 ;
        RECT 13.415 -0.085 13.585 0.085 ;
        RECT 13.775 -0.085 13.945 0.085 ;
        RECT 14.135 -0.085 14.305 0.085 ;
        RECT 14.495 -0.085 14.665 0.085 ;
        RECT 14.855 -0.085 15.025 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 15.120 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 15.120 6.205 ;
        RECT 9.915 5.200 10.085 6.035 ;
        RECT 12.075 5.200 12.245 6.035 ;
        RECT 9.835 5.030 10.165 5.200 ;
        RECT 11.995 5.030 12.325 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
        RECT 10.895 6.035 11.065 6.205 ;
        RECT 11.255 6.035 11.425 6.205 ;
        RECT 11.615 6.035 11.785 6.205 ;
        RECT 11.975 6.035 12.145 6.205 ;
        RECT 12.335 6.035 12.505 6.205 ;
        RECT 12.695 6.035 12.865 6.205 ;
        RECT 13.055 6.035 13.225 6.205 ;
        RECT 13.415 6.035 13.585 6.205 ;
        RECT 13.775 6.035 13.945 6.205 ;
        RECT 14.135 6.035 14.305 6.205 ;
        RECT 14.495 6.035 14.665 6.205 ;
        RECT 14.855 6.035 15.025 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 15.120 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 15.300 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 5.955 1.445 ;
      LAYER li1 ;
        RECT 2.275 5.030 8.465 5.200 ;
        RECT 0.115 4.690 3.685 4.860 ;
        RECT 8.295 4.390 8.465 5.030 ;
        RECT 8.755 4.690 14.485 4.860 ;
        RECT 5.515 4.220 6.925 4.390 ;
        RECT 7.675 4.220 8.005 4.390 ;
        RECT 8.295 4.220 11.245 4.390 ;
        RECT 13.075 4.220 13.405 4.390 ;
        RECT 7.755 3.230 7.925 4.220 ;
        RECT 13.155 3.230 13.325 4.220 ;
        RECT 7.755 3.060 13.325 3.230 ;
  END
END NR4D1_2

#--------EOF---------

MACRO NR4D1_3
  CLASS CORE ;
  FOREIGN NR4D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.040 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.869300 ;
    PORT
      LAYER li1 ;
        RECT 1.275 4.220 3.685 4.390 ;
        RECT 1.275 1.500 1.445 4.220 ;
        RECT 1.275 1.330 3.605 1.500 ;
        RECT 1.275 1.090 1.445 1.330 ;
        RECT 3.435 1.090 3.605 1.330 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END zn
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 0.735 0.440 0.905 1.090 ;
        RECT 0.655 0.270 0.985 0.440 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 1.735 1.980 12.865 2.150 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 2.815 3.060 6.385 3.230 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.398250 ;
    PORT
      LAYER li1 ;
        RECT 3.895 2.520 4.685 2.690 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 14.040 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
        RECT 8.735 -0.085 8.905 0.085 ;
        RECT 9.095 -0.085 9.265 0.085 ;
        RECT 9.455 -0.085 9.625 0.085 ;
        RECT 9.815 -0.085 9.985 0.085 ;
        RECT 10.175 -0.085 10.345 0.085 ;
        RECT 10.535 -0.085 10.705 0.085 ;
        RECT 10.895 -0.085 11.065 0.085 ;
        RECT 11.255 -0.085 11.425 0.085 ;
        RECT 11.615 -0.085 11.785 0.085 ;
        RECT 11.975 -0.085 12.145 0.085 ;
        RECT 12.335 -0.085 12.505 0.085 ;
        RECT 12.695 -0.085 12.865 0.085 ;
        RECT 13.055 -0.085 13.225 0.085 ;
        RECT 13.415 -0.085 13.585 0.085 ;
        RECT 13.775 -0.085 13.945 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 14.040 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 14.040 6.205 ;
        RECT 8.835 5.200 9.005 6.035 ;
        RECT 10.995 5.200 11.165 6.035 ;
        RECT 8.755 5.030 9.085 5.200 ;
        RECT 10.915 5.030 11.245 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
        RECT 8.735 6.035 8.905 6.205 ;
        RECT 9.095 6.035 9.265 6.205 ;
        RECT 9.455 6.035 9.625 6.205 ;
        RECT 9.815 6.035 9.985 6.205 ;
        RECT 10.175 6.035 10.345 6.205 ;
        RECT 10.535 6.035 10.705 6.205 ;
        RECT 10.895 6.035 11.065 6.205 ;
        RECT 11.255 6.035 11.425 6.205 ;
        RECT 11.615 6.035 11.785 6.205 ;
        RECT 11.975 6.035 12.145 6.205 ;
        RECT 12.335 6.035 12.505 6.205 ;
        RECT 12.695 6.035 12.865 6.205 ;
        RECT 13.055 6.035 13.225 6.205 ;
        RECT 13.415 6.035 13.585 6.205 ;
        RECT 13.775 6.035 13.945 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 14.040 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 14.220 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 4.875 1.445 ;
      LAYER li1 ;
        RECT 0.115 4.690 10.165 4.860 ;
        RECT 11.535 4.690 13.405 4.860 ;
        RECT 11.535 4.390 11.705 4.690 ;
        RECT 4.435 4.220 5.845 4.390 ;
        RECT 6.595 4.220 6.925 4.390 ;
        RECT 7.675 4.220 11.705 4.390 ;
        RECT 11.995 4.220 12.325 4.390 ;
        RECT 6.675 3.230 6.845 4.220 ;
        RECT 12.075 3.230 12.245 4.220 ;
        RECT 6.675 3.060 12.245 3.230 ;
  END
END NR4D1_3

#--------EOF---------

MACRO OA21D1
  CLASS CORE ;
  FOREIGN OA21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.815 2.520 3.605 2.690 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 4.435 4.220 4.765 4.390 ;
        RECT 4.515 1.090 4.685 4.220 ;
        RECT 4.435 0.920 4.765 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 0.000 -0.085 6.480 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.480 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 6.480 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 6.480 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 6.660 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 5.955 1.690 ;
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 1.275 3.230 1.445 4.220 ;
        RECT 1.275 3.060 4.225 3.230 ;
        RECT 2.355 2.150 2.525 3.060 ;
        RECT 2.355 1.980 3.685 2.150 ;
        RECT 2.355 1.090 2.525 1.980 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 1.275 0.440 1.445 0.920 ;
        RECT 3.435 0.440 3.605 0.920 ;
        RECT 1.275 0.270 3.605 0.440 ;
  END
END OA21D1

#--------EOF---------

MACRO OA21D1_1
  CLASS CORE ;
  FOREIGN OA21D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 4.435 4.220 4.765 4.390 ;
        RECT 4.515 1.090 4.685 4.220 ;
        RECT 4.435 0.920 4.765 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 0.000 -0.085 6.480 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.480 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 6.480 6.205 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 6.480 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 6.660 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 5.955 1.690 ;
      LAYER li1 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 0.195 3.230 0.365 4.220 ;
        RECT 3.435 3.230 3.605 4.220 ;
        RECT 0.195 3.060 3.685 3.230 ;
        RECT 1.275 1.090 1.445 3.060 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 0.195 0.440 0.365 0.920 ;
        RECT 2.355 0.440 2.525 0.920 ;
        RECT 0.195 0.270 2.525 0.440 ;
  END
END OA21D1_1

#--------EOF---------

MACRO OA21D1_2
  CLASS CORE ;
  FOREIGN OA21D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 3.975 2.150 4.145 2.690 ;
        RECT 3.895 1.980 4.225 2.150 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 5.515 4.220 5.845 4.390 ;
        RECT 5.595 1.090 5.765 4.220 ;
        RECT 5.515 0.920 5.845 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 6.480 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.480 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 6.480 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 6.480 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 6.660 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 5.955 1.690 ;
      LAYER li1 ;
        RECT 2.275 4.220 3.685 4.390 ;
        RECT 1.275 1.330 3.605 1.500 ;
        RECT 1.275 1.090 1.445 1.330 ;
        RECT 3.435 1.090 3.605 1.330 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 0.195 0.440 0.365 0.920 ;
        RECT 2.355 0.440 2.525 0.920 ;
        RECT 0.115 0.270 0.445 0.440 ;
        RECT 2.275 0.270 2.605 0.440 ;
  END
END OA21D1_2

#--------EOF---------

MACRO OA21D1_3
  CLASS CORE ;
  FOREIGN OA21D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.480 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 4.435 4.220 4.765 4.390 ;
        RECT 4.515 1.090 4.685 4.220 ;
        RECT 4.435 0.920 4.765 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 5.595 0.085 5.765 0.920 ;
        RECT 0.000 -0.085 6.480 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.480 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 6.480 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 5.595 5.200 5.765 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 6.480 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 6.660 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 5.955 1.690 ;
      LAYER li1 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 0.195 3.230 0.365 4.220 ;
        RECT 3.435 3.230 3.605 4.220 ;
        RECT 0.195 3.060 3.685 3.230 ;
        RECT 2.355 1.090 2.525 3.060 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 1.275 0.440 1.445 0.920 ;
        RECT 3.435 0.440 3.605 0.920 ;
        RECT 1.275 0.270 3.605 0.440 ;
  END
END OA21D1_3

#--------EOF---------

MACRO OAI21D1
  CLASS CORE ;
  FOREIGN OAI21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.674000 ;
    PORT
      LAYER li1 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 1.275 3.230 1.445 4.220 ;
        RECT 1.275 3.060 2.525 3.230 ;
        RECT 2.355 1.090 2.525 3.060 ;
        RECT 2.275 0.920 2.605 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.320 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 4.320 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 3.355 5.030 3.685 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 4.320 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 4.500 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 3.795 1.690 ;
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 1.275 0.440 1.445 0.920 ;
        RECT 3.435 0.440 3.605 0.920 ;
        RECT 1.275 0.270 3.605 0.440 ;
  END
END OAI21D1

#--------EOF---------

MACRO OAI21D1_1
  CLASS CORE ;
  FOREIGN OAI21D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.674000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 4.220 2.605 4.390 ;
        RECT 2.355 2.150 2.525 4.220 ;
        RECT 1.275 1.980 2.525 2.150 ;
        RECT 1.275 1.090 1.445 1.980 ;
        RECT 1.195 0.920 1.525 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.690 1.985 3.230 ;
        RECT 1.735 2.520 2.065 2.690 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.320 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 4.320 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 3.355 5.030 3.685 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 4.320 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 4.500 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 3.795 1.690 ;
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 0.195 0.440 0.365 0.920 ;
        RECT 2.355 0.440 2.525 0.920 ;
        RECT 0.195 0.270 2.525 0.440 ;
  END
END OAI21D1_1

#--------EOF---------

MACRO OAI21D1_2
  CLASS CORE ;
  FOREIGN OAI21D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.196000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 4.220 3.685 4.390 ;
        RECT 0.195 1.090 0.365 4.220 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 0.195 0.440 0.365 0.920 ;
        RECT 2.355 0.440 2.525 0.920 ;
        RECT 0.195 0.270 2.525 0.440 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 3.975 2.150 4.145 2.690 ;
        RECT 3.895 1.980 4.225 2.150 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 5.400 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.400 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 5.400 6.205 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 5.400 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 5.580 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 4.875 1.690 ;
      LAYER li1 ;
        RECT 1.275 1.330 3.605 1.500 ;
        RECT 1.275 1.090 1.445 1.330 ;
        RECT 3.435 1.090 3.605 1.330 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
  END
END OAI21D1_2

#--------EOF---------

MACRO OAI21D1_3
  CLASS CORE ;
  FOREIGN OAI21D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.196000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 4.220 3.685 4.390 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 3.145 1.090 ;
        RECT 0.195 0.440 0.365 0.920 ;
        RECT 2.355 0.440 2.525 0.920 ;
        RECT 0.195 0.270 2.525 0.440 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 3.975 2.150 4.145 2.690 ;
        RECT 3.895 1.980 4.225 2.150 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 5.400 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.400 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 5.400 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 5.400 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 5.580 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 4.875 1.690 ;
      LAYER li1 ;
        RECT 1.275 1.330 3.605 1.500 ;
        RECT 1.275 1.090 1.445 1.330 ;
        RECT 3.435 1.090 3.605 1.330 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
  END
END OAI21D1_3

#--------EOF---------

MACRO OR2D1
  CLASS CORE ;
  FOREIGN OR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.058350 ;
    PORT
      LAYER li1 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 3.435 1.090 3.605 4.220 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 0.000 -0.085 4.320 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.320 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 4.320 6.205 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 2.275 5.030 2.605 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 4.320 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 4.500 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 3.795 1.625 ;
      LAYER li1 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 0.195 3.230 0.365 4.220 ;
        RECT 0.195 3.060 3.145 3.230 ;
        RECT 1.275 1.090 1.445 3.060 ;
        RECT 1.195 0.920 1.525 1.090 ;
  END
END OR2D1

#--------EOF---------

MACRO OR2D1_1
  CLASS CORE ;
  FOREIGN OR2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.058350 ;
    PORT
      LAYER li1 ;
        RECT 3.355 4.220 4.145 4.390 ;
        RECT 3.975 1.090 4.145 4.220 ;
        RECT 3.355 0.920 4.145 1.090 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 2.355 0.085 2.525 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 5.400 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.400 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 5.400 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 5.400 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 5.580 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 4.875 1.625 ;
      LAYER li1 ;
        RECT 2.275 4.220 2.605 4.390 ;
        RECT 2.355 3.230 2.525 4.220 ;
        RECT 1.275 3.060 3.685 3.230 ;
        RECT 1.275 1.090 1.445 3.060 ;
        RECT 1.195 0.920 1.525 1.090 ;
  END
END OR2D1_1

#--------EOF---------

MACRO OR2D1_2
  CLASS CORE ;
  FOREIGN OR2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.058350 ;
    PORT
      LAYER li1 ;
        RECT 2.815 4.220 3.685 4.390 ;
        RECT 2.815 0.920 3.685 1.090 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.690 0.905 3.230 ;
        RECT 0.655 2.520 0.985 2.690 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.690 1.985 3.230 ;
        RECT 1.735 2.520 2.065 2.690 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 5.400 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.400 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 5.400 6.205 ;
        RECT 2.355 5.200 2.525 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 5.400 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 5.580 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 4.875 1.625 ;
      LAYER li1 ;
        RECT 0.115 4.220 2.525 4.390 ;
        RECT 2.355 2.150 2.525 4.220 ;
        RECT 0.195 1.980 4.225 2.150 ;
        RECT 0.195 1.090 0.365 1.980 ;
        RECT 2.355 1.090 2.525 1.980 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 2.355 0.440 2.525 0.920 ;
        RECT 2.355 0.270 4.225 0.440 ;
  END
END OR2D1_2

#--------EOF---------

MACRO OR2D1_3
  CLASS CORE ;
  FOREIGN OR2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.400 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.058350 ;
    PORT
      LAYER li1 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 3.435 1.090 3.605 4.220 ;
        RECT 3.355 0.920 3.685 1.090 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.150 1.985 2.690 ;
        RECT 1.735 1.980 2.065 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.260250 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 0.000 -0.085 5.400 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.400 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 5.400 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 5.400 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 5.580 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 4.875 1.625 ;
      LAYER li1 ;
        RECT 2.275 4.220 2.605 4.390 ;
        RECT 2.355 3.230 2.525 4.220 ;
        RECT 2.275 3.060 2.605 3.230 ;
        RECT 2.355 1.500 2.525 3.060 ;
        RECT 0.195 1.330 2.525 1.500 ;
        RECT 0.195 1.090 0.365 1.330 ;
        RECT 2.355 1.090 2.525 1.330 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
  END
END OR2D1_3

#--------EOF---------

MACRO TIEH
  CLASS CORE ;
  FOREIGN TIEH ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.160 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.195 4.220 0.365 5.200 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 0.000 -0.085 2.160 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 2.160 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 2.160 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 2.160 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 2.340 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 1.635 1.690 ;
      LAYER li1 ;
        RECT 0.115 0.920 0.905 1.090 ;
        RECT 0.735 0.440 0.905 0.920 ;
        RECT 0.655 0.270 0.985 0.440 ;
  END
END TIEH

#--------EOF---------

MACRO TIEL
  CLASS CORE ;
  FOREIGN TIEL ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.160 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.090 0.905 1.500 ;
        RECT 0.195 0.920 0.905 1.090 ;
    END
  END zn
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 1.275 0.085 1.445 0.920 ;
        RECT 0.000 -0.085 2.160 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 2.160 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 2.160 6.205 ;
        RECT 1.275 5.200 1.445 6.035 ;
        RECT 1.195 5.030 1.525 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 2.160 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 2.340 6.445 ;
      LAYER pwell ;
        RECT 0.005 0.730 1.635 1.690 ;
      LAYER li1 ;
        RECT 0.115 4.220 0.445 4.390 ;
        RECT 0.195 3.230 0.365 4.220 ;
        RECT 0.115 3.060 0.445 3.230 ;
  END
END TIEL

#--------EOF---------

MACRO XNR2D1
  CLASS CORE ;
  FOREIGN XNR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 6.595 4.220 6.925 4.390 ;
        RECT 6.675 1.090 6.845 4.220 ;
        RECT 6.595 0.920 6.925 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.291000 ;
    PORT
      LAYER li1 ;
        RECT 4.975 4.220 5.305 4.390 ;
        RECT 5.055 2.690 5.225 4.220 ;
        RECT 4.975 2.520 5.305 2.690 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 7.675 0.920 8.005 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 7.755 0.085 7.925 0.920 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.640 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 8.640 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 7.755 5.200 7.925 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 8.640 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 8.820 6.445 ;
      LAYER pwell ;
        RECT 0.005 1.410 1.635 1.690 ;
        RECT 6.485 1.410 8.115 1.690 ;
        RECT 0.005 0.730 8.115 1.410 ;
      LAYER li1 ;
        RECT 2.275 5.030 3.065 5.200 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 1.195 4.220 2.605 4.390 ;
        RECT 1.275 1.090 1.445 4.220 ;
        RECT 2.895 3.230 3.065 5.030 ;
        RECT 2.355 3.060 3.145 3.230 ;
        RECT 2.355 1.090 2.525 3.060 ;
        RECT 3.435 2.690 3.605 5.030 ;
        RECT 3.895 4.220 4.225 4.390 ;
        RECT 3.975 2.690 4.145 4.220 ;
        RECT 2.895 2.520 3.605 2.690 ;
        RECT 3.895 2.520 4.225 2.690 ;
        RECT 2.895 1.090 3.065 2.520 ;
        RECT 5.595 2.150 5.765 5.030 ;
        RECT 3.355 1.980 5.765 2.150 ;
        RECT 5.595 1.090 5.765 1.980 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 2.895 0.920 3.685 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
  END
END XNR2D1

#--------EOF---------

MACRO XNR2D1_1
  CLASS CORE ;
  FOREIGN XNR2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 3.975 3.230 4.145 4.390 ;
        RECT 3.895 3.060 4.225 3.230 ;
    END
  END a2
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 6.595 4.220 6.925 4.390 ;
        RECT 6.675 1.090 6.845 4.220 ;
        RECT 6.595 0.920 6.925 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.291000 ;
    PORT
      LAYER li1 ;
        RECT 1.735 5.680 2.065 5.850 ;
        RECT 1.815 4.860 1.985 5.680 ;
        RECT 1.815 4.690 5.225 4.860 ;
        RECT 5.055 4.390 5.225 4.690 ;
        RECT 4.975 4.220 5.305 4.390 ;
        RECT 2.815 1.980 5.305 2.150 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 7.675 0.920 8.005 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 7.755 0.085 7.925 0.920 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.640 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 8.640 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 7.755 5.200 7.925 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 8.640 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 8.820 6.445 ;
      LAYER pwell ;
        RECT 3.245 1.410 4.875 1.690 ;
        RECT 6.485 1.410 8.115 1.690 ;
        RECT 0.005 0.730 8.115 1.410 ;
      LAYER li1 ;
        RECT 2.275 5.680 2.605 5.850 ;
        RECT 2.355 5.200 2.525 5.680 ;
        RECT 0.735 5.030 1.525 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 0.735 1.090 0.905 5.030 ;
        RECT 3.355 4.220 3.685 4.390 ;
        RECT 3.435 3.230 3.605 4.220 ;
        RECT 1.195 3.060 3.605 3.230 ;
        RECT 5.595 2.690 5.765 5.030 ;
        RECT 2.815 2.520 5.765 2.690 ;
        RECT 1.815 1.330 3.605 1.500 ;
        RECT 0.735 0.920 1.525 1.090 ;
        RECT 1.815 0.440 1.985 1.330 ;
        RECT 3.435 1.090 3.605 1.330 ;
        RECT 5.595 1.090 5.765 2.520 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 2.355 0.440 2.525 0.920 ;
        RECT 0.655 0.270 1.985 0.440 ;
        RECT 2.275 0.270 2.605 0.440 ;
  END
END XNR2D1_1

#--------EOF---------

MACRO XNR2D1_2
  CLASS CORE ;
  FOREIGN XNR2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 3.435 2.690 3.605 3.230 ;
        RECT 3.355 2.520 3.685 2.690 ;
    END
  END a2
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 7.675 4.220 8.005 4.390 ;
        RECT 7.755 1.090 7.925 4.220 ;
        RECT 7.675 0.920 8.005 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.291000 ;
    PORT
      LAYER li1 ;
        RECT 3.975 0.440 4.145 1.090 ;
        RECT 3.895 0.270 4.225 0.440 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 6.595 0.920 6.925 1.090 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 6.675 0.085 6.845 0.920 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.640 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 8.640 6.205 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 6.675 5.200 6.845 6.035 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 6.595 5.030 6.925 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 8.640 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 8.820 6.445 ;
      LAYER pwell ;
        RECT 2.165 1.410 3.795 1.690 ;
        RECT 6.485 1.410 8.115 1.690 ;
        RECT 0.005 0.730 8.115 1.410 ;
      LAYER li1 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 0.195 4.860 0.365 5.030 ;
        RECT 5.595 4.860 5.765 5.030 ;
        RECT 0.195 4.690 5.765 4.860 ;
        RECT 0.735 1.090 0.905 4.690 ;
        RECT 2.275 4.220 2.605 4.390 ;
        RECT 2.355 1.090 2.525 4.220 ;
        RECT 2.895 2.150 3.065 4.690 ;
        RECT 2.895 1.980 4.765 2.150 ;
        RECT 2.895 1.330 6.305 1.500 ;
        RECT 2.895 1.090 3.065 1.330 ;
        RECT 0.115 0.920 0.905 1.090 ;
        RECT 2.275 0.920 3.065 1.090 ;
        RECT 4.975 0.920 5.845 1.090 ;
        RECT 6.135 0.440 6.305 1.330 ;
        RECT 6.055 0.270 6.385 0.440 ;
  END
END XNR2D1_2

#--------EOF---------

MACRO XNR2D1_3
  CLASS CORE ;
  FOREIGN XNR2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.150 3.065 2.690 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END a2
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 5.515 4.220 5.845 4.390 ;
        RECT 5.595 1.090 5.765 4.220 ;
        RECT 5.515 0.920 5.845 1.090 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.291000 ;
    PORT
      LAYER li1 ;
        RECT 3.975 0.440 4.145 1.090 ;
        RECT 3.895 0.270 4.225 0.440 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 6.595 0.920 6.925 1.090 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 6.675 0.085 6.845 0.920 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.640 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 8.640 6.205 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 6.675 5.200 6.845 6.035 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 6.595 5.030 6.925 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 8.640 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 8.820 6.445 ;
      LAYER pwell ;
        RECT 2.165 1.410 3.795 1.690 ;
        RECT 5.405 1.410 7.035 1.690 ;
        RECT 0.005 0.730 8.115 1.410 ;
      LAYER li1 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
        RECT 0.195 4.860 0.365 5.030 ;
        RECT 7.755 4.860 7.925 5.030 ;
        RECT 0.195 4.690 7.925 4.860 ;
        RECT 1.815 2.150 1.985 4.690 ;
        RECT 2.275 4.220 2.605 4.390 ;
        RECT 0.735 1.980 1.985 2.150 ;
        RECT 0.735 1.090 0.905 1.980 ;
        RECT 2.355 1.090 2.525 4.220 ;
        RECT 6.135 1.500 6.305 4.690 ;
        RECT 2.895 1.330 5.225 1.500 ;
        RECT 6.135 1.330 7.385 1.500 ;
        RECT 2.895 1.090 3.065 1.330 ;
        RECT 0.115 0.920 0.905 1.090 ;
        RECT 2.275 0.920 3.065 1.090 ;
        RECT 5.055 0.440 5.225 1.330 ;
        RECT 7.215 1.090 7.385 1.330 ;
        RECT 7.215 0.920 8.005 1.090 ;
        RECT 5.055 0.270 6.385 0.440 ;
  END
END XNR2D1_3

#--------EOF---------

MACRO XOR2D1
  CLASS CORE ;
  FOREIGN XOR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.291000 ;
    PORT
      LAYER li1 ;
        RECT 2.815 2.520 5.305 2.690 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 6.595 4.220 6.925 4.390 ;
        RECT 6.675 1.090 6.845 4.220 ;
        RECT 6.595 0.920 6.925 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 7.675 0.920 8.005 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 7.755 0.085 7.925 0.920 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.640 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 8.640 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 7.755 5.200 7.925 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 8.640 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 8.820 6.445 ;
      LAYER pwell ;
        RECT 3.245 1.410 4.875 1.690 ;
        RECT 6.485 1.410 8.115 1.690 ;
        RECT 0.005 0.730 8.115 1.410 ;
      LAYER li1 ;
        RECT 0.655 5.680 3.605 5.850 ;
        RECT 3.435 5.200 3.605 5.680 ;
        RECT 1.195 5.030 1.525 5.200 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 1.275 1.090 1.445 5.030 ;
        RECT 1.735 4.220 2.065 4.390 ;
        RECT 1.815 2.150 1.985 4.220 ;
        RECT 2.355 3.230 2.525 5.030 ;
        RECT 2.355 3.060 5.305 3.230 ;
        RECT 5.595 2.150 5.765 5.030 ;
        RECT 1.815 1.980 5.765 2.150 ;
        RECT 2.355 1.330 6.305 1.500 ;
        RECT 2.355 1.090 2.525 1.330 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 3.435 0.440 3.605 0.920 ;
        RECT 5.595 0.440 5.765 0.920 ;
        RECT 6.135 0.440 6.305 1.330 ;
        RECT 0.655 0.270 3.605 0.440 ;
        RECT 5.515 0.270 5.845 0.440 ;
        RECT 6.055 0.270 6.385 0.440 ;
  END
END XOR2D1

#--------EOF---------

MACRO XOR2D1_1
  CLASS CORE ;
  FOREIGN XOR2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.291000 ;
    PORT
      LAYER li1 ;
        RECT 0.655 0.270 1.445 0.440 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 3.230 3.065 4.390 ;
        RECT 2.815 3.060 3.145 3.230 ;
    END
  END a2
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 7.675 4.220 8.005 4.390 ;
        RECT 7.755 1.090 7.925 4.220 ;
        RECT 7.675 0.920 8.005 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 6.595 0.920 6.925 1.090 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 6.675 0.085 6.845 0.920 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.640 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 8.640 6.205 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 6.675 5.200 6.845 6.035 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 6.595 5.030 6.925 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 8.640 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 8.820 6.445 ;
      LAYER pwell ;
        RECT 2.165 1.410 3.795 1.690 ;
        RECT 6.485 1.410 8.115 1.690 ;
        RECT 0.005 0.730 8.115 1.410 ;
      LAYER li1 ;
        RECT 0.655 5.680 1.985 5.850 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 1.195 5.030 1.525 5.200 ;
        RECT 0.195 1.090 0.365 5.030 ;
        RECT 1.275 1.500 1.445 5.030 ;
        RECT 1.815 3.230 1.985 5.680 ;
        RECT 4.435 5.030 4.765 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 1.735 3.060 2.065 3.230 ;
        RECT 4.515 2.690 4.685 5.030 ;
        RECT 2.275 2.520 5.305 2.690 ;
        RECT 2.355 1.980 5.305 2.150 ;
        RECT 2.355 1.500 2.525 1.980 ;
        RECT 5.595 1.500 5.765 5.030 ;
        RECT 6.055 2.520 6.385 2.690 ;
        RECT 1.275 1.330 2.525 1.500 ;
        RECT 2.895 1.330 5.765 1.500 ;
        RECT 1.275 1.090 1.445 1.330 ;
        RECT 2.895 1.090 3.065 1.330 ;
        RECT 5.595 1.090 5.765 1.330 ;
        RECT 0.115 0.920 3.065 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 4.515 0.440 4.685 0.920 ;
        RECT 6.135 0.440 6.305 2.520 ;
        RECT 4.515 0.270 6.305 0.440 ;
  END
END XOR2D1_1

#--------EOF---------

MACRO XOR2D1_2
  CLASS CORE ;
  FOREIGN XOR2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.291000 ;
    PORT
      LAYER li1 ;
        RECT 0.655 0.270 1.445 0.440 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.690 3.065 3.230 ;
        RECT 2.815 2.520 3.145 2.690 ;
    END
  END a2
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 5.515 4.220 5.845 4.390 ;
        RECT 5.595 1.090 5.765 4.220 ;
        RECT 5.515 0.920 5.845 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 6.595 0.920 6.925 1.090 ;
        RECT 3.435 0.085 3.605 0.920 ;
        RECT 6.675 0.085 6.845 0.920 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.640 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 8.640 6.205 ;
        RECT 3.435 5.200 3.605 6.035 ;
        RECT 6.675 5.200 6.845 6.035 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 6.595 5.030 6.925 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 8.640 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 8.820 6.445 ;
      LAYER pwell ;
        RECT 2.165 1.410 3.795 1.690 ;
        RECT 5.405 1.410 7.035 1.690 ;
        RECT 0.005 0.730 8.115 1.410 ;
      LAYER li1 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 1.195 5.030 1.525 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
        RECT 0.195 1.090 0.365 5.030 ;
        RECT 1.275 1.500 1.445 5.030 ;
        RECT 2.355 1.980 5.305 2.150 ;
        RECT 2.355 1.500 2.525 1.980 ;
        RECT 1.275 1.330 2.525 1.500 ;
        RECT 2.895 1.330 5.225 1.500 ;
        RECT 1.275 1.090 1.445 1.330 ;
        RECT 2.895 1.090 3.065 1.330 ;
        RECT 0.115 0.920 3.065 1.090 ;
        RECT 5.055 0.440 5.225 1.330 ;
        RECT 7.755 1.090 7.925 5.030 ;
        RECT 7.675 0.920 8.005 1.090 ;
        RECT 7.755 0.440 7.925 0.920 ;
        RECT 5.055 0.270 6.385 0.440 ;
        RECT 7.675 0.270 8.005 0.440 ;
  END
END XOR2D1_2

#--------EOF---------

MACRO XOR2D1_3
  CLASS CORE ;
  FOREIGN XOR2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 6.120 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.291000 ;
    PORT
      LAYER li1 ;
        RECT 2.815 5.680 3.145 5.850 ;
        RECT 2.895 2.150 3.065 5.680 ;
        RECT 2.815 1.980 3.145 2.150 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.150 0.905 2.690 ;
        RECT 0.655 1.980 0.985 2.150 ;
    END
  END a2
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.098000 ;
    PORT
      LAYER li1 ;
        RECT 6.595 4.220 6.925 4.390 ;
        RECT 6.675 1.090 6.845 4.220 ;
        RECT 6.595 0.920 6.925 1.090 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.920 0.445 1.090 ;
        RECT 4.435 0.920 4.765 1.090 ;
        RECT 7.675 0.920 8.005 1.090 ;
        RECT 0.195 0.085 0.365 0.920 ;
        RECT 4.515 0.085 4.685 0.920 ;
        RECT 7.755 0.085 7.925 0.920 ;
        RECT 0.000 -0.085 8.640 0.085 ;
      LAYER mcon ;
        RECT 0.095 -0.085 0.265 0.085 ;
        RECT 0.455 -0.085 0.625 0.085 ;
        RECT 0.815 -0.085 0.985 0.085 ;
        RECT 1.175 -0.085 1.345 0.085 ;
        RECT 1.535 -0.085 1.705 0.085 ;
        RECT 1.895 -0.085 2.065 0.085 ;
        RECT 2.255 -0.085 2.425 0.085 ;
        RECT 2.615 -0.085 2.785 0.085 ;
        RECT 2.975 -0.085 3.145 0.085 ;
        RECT 3.335 -0.085 3.505 0.085 ;
        RECT 3.695 -0.085 3.865 0.085 ;
        RECT 4.055 -0.085 4.225 0.085 ;
        RECT 4.415 -0.085 4.585 0.085 ;
        RECT 4.775 -0.085 4.945 0.085 ;
        RECT 5.135 -0.085 5.305 0.085 ;
        RECT 5.495 -0.085 5.665 0.085 ;
        RECT 5.855 -0.085 6.025 0.085 ;
        RECT 6.215 -0.085 6.385 0.085 ;
        RECT 6.575 -0.085 6.745 0.085 ;
        RECT 6.935 -0.085 7.105 0.085 ;
        RECT 7.295 -0.085 7.465 0.085 ;
        RECT 7.655 -0.085 7.825 0.085 ;
        RECT 8.015 -0.085 8.185 0.085 ;
        RECT 8.375 -0.085 8.545 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.640 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 6.035 8.640 6.205 ;
        RECT 0.195 5.200 0.365 6.035 ;
        RECT 4.515 5.200 4.685 6.035 ;
        RECT 7.755 5.200 7.925 6.035 ;
        RECT 0.115 5.030 0.445 5.200 ;
        RECT 4.435 5.030 4.765 5.200 ;
        RECT 7.675 5.030 8.005 5.200 ;
      LAYER mcon ;
        RECT 0.095 6.035 0.265 6.205 ;
        RECT 0.455 6.035 0.625 6.205 ;
        RECT 0.815 6.035 0.985 6.205 ;
        RECT 1.175 6.035 1.345 6.205 ;
        RECT 1.535 6.035 1.705 6.205 ;
        RECT 1.895 6.035 2.065 6.205 ;
        RECT 2.255 6.035 2.425 6.205 ;
        RECT 2.615 6.035 2.785 6.205 ;
        RECT 2.975 6.035 3.145 6.205 ;
        RECT 3.335 6.035 3.505 6.205 ;
        RECT 3.695 6.035 3.865 6.205 ;
        RECT 4.055 6.035 4.225 6.205 ;
        RECT 4.415 6.035 4.585 6.205 ;
        RECT 4.775 6.035 4.945 6.205 ;
        RECT 5.135 6.035 5.305 6.205 ;
        RECT 5.495 6.035 5.665 6.205 ;
        RECT 5.855 6.035 6.025 6.205 ;
        RECT 6.215 6.035 6.385 6.205 ;
        RECT 6.575 6.035 6.745 6.205 ;
        RECT 6.935 6.035 7.105 6.205 ;
        RECT 7.295 6.035 7.465 6.205 ;
        RECT 7.655 6.035 7.825 6.205 ;
        RECT 8.015 6.035 8.185 6.205 ;
        RECT 8.375 6.035 8.545 6.205 ;
      LAYER met1 ;
        RECT 0.000 5.985 8.640 6.255 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 2.860 8.820 6.445 ;
      LAYER pwell ;
        RECT 0.005 1.410 1.635 1.690 ;
        RECT 6.485 1.410 8.115 1.690 ;
        RECT 0.005 0.730 8.115 1.410 ;
      LAYER li1 ;
        RECT 2.275 5.030 2.605 5.200 ;
        RECT 3.355 5.030 3.685 5.200 ;
        RECT 5.515 5.030 5.845 5.200 ;
        RECT 1.195 4.220 1.525 4.390 ;
        RECT 1.275 2.690 1.445 4.220 ;
        RECT 1.275 2.520 2.065 2.690 ;
        RECT 1.275 1.090 1.445 2.520 ;
        RECT 2.355 1.090 2.525 5.030 ;
        RECT 3.435 1.090 3.605 5.030 ;
        RECT 3.895 4.220 4.225 4.390 ;
        RECT 3.975 2.690 4.145 4.220 ;
        RECT 5.595 3.230 5.765 5.030 ;
        RECT 4.435 3.060 5.765 3.230 ;
        RECT 3.895 2.520 4.225 2.690 ;
        RECT 5.595 1.090 5.765 3.060 ;
        RECT 1.195 0.920 1.525 1.090 ;
        RECT 2.275 0.920 2.605 1.090 ;
        RECT 3.355 0.920 3.685 1.090 ;
        RECT 5.515 0.920 5.845 1.090 ;
        RECT 2.355 0.440 2.525 0.920 ;
        RECT 2.275 0.270 2.605 0.440 ;
  END
END XOR2D1_3

#--------EOF---------


END LIBRARY
