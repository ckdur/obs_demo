VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

SITE obssite
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.34 BY 4.08 ;
END obssite

#--------EOF---------

MACRO AN2D1
  CLASS CORE ;
  FOREIGN AN2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 3.355 2.545 3.685 2.715 ;
        RECT 3.435 1.185 3.605 2.545 ;
        RECT 3.355 1.015 3.685 1.185 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 0.000 -0.085 5.440 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 5.440 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 5.440 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 5.620 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.545 4.875 1.395 ;
        RECT 3.245 0.485 4.875 0.545 ;
      LAYER li1 ;
        RECT 1.195 2.545 2.525 2.715 ;
        RECT 2.355 1.765 2.525 2.545 ;
        RECT 2.275 1.595 2.605 1.765 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 2.275 1.015 2.605 1.185 ;
  END
END AN2D1

#--------EOF---------

MACRO AN2D1_1
  CLASS CORE ;
  FOREIGN AN2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.080 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.002000 ;
    PORT
      LAYER li1 ;
        RECT 3.355 2.545 3.685 2.715 ;
        RECT 3.435 1.185 3.605 2.545 ;
        RECT 3.355 1.015 3.685 1.185 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 0.000 -0.085 4.080 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.080 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 4.080 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 2.275 2.885 2.605 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 4.080 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 4.260 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.545 3.795 1.395 ;
        RECT 2.165 0.485 3.795 0.545 ;
      LAYER li1 ;
        RECT 1.195 2.545 3.065 2.715 ;
        RECT 1.275 2.445 1.445 2.545 ;
        RECT 2.895 2.445 3.065 2.545 ;
        RECT 0.195 2.275 1.445 2.445 ;
        RECT 2.815 2.275 3.145 2.445 ;
        RECT 0.195 1.185 0.365 2.275 ;
        RECT 0.115 1.015 0.445 1.185 ;
  END
END AN2D1_1

#--------EOF---------

MACRO AN2D1_2
  CLASS CORE ;
  FOREIGN AN2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 3.355 2.545 3.685 2.715 ;
        RECT 3.435 1.185 3.605 2.545 ;
        RECT 3.355 1.015 3.685 1.185 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.105 0.905 2.445 ;
        RECT 0.655 1.935 0.985 2.105 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 0.000 -0.085 5.440 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 5.440 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 5.440 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 5.620 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.545 4.875 1.395 ;
        RECT 3.245 0.485 4.875 0.545 ;
      LAYER li1 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 2.275 2.545 2.605 2.715 ;
        RECT 0.195 1.765 0.365 2.545 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 2.275 2.275 2.605 2.445 ;
        RECT 2.355 1.765 2.525 2.275 ;
        RECT 0.195 1.595 3.145 1.765 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 2.275 1.015 2.605 1.185 ;
  END
END AN2D1_2

#--------EOF---------

MACRO AN2D1_3
  CLASS CORE ;
  FOREIGN AN2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 3.355 2.545 3.685 2.715 ;
        RECT 3.435 1.185 3.605 2.545 ;
        RECT 3.355 1.015 3.685 1.185 ;
    END
  END z
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.935 2.605 2.105 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 0.000 -0.085 5.440 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 5.440 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 5.440 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 5.620 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.545 4.875 1.395 ;
        RECT 3.245 0.485 4.875 0.545 ;
      LAYER li1 ;
        RECT 0.115 2.545 1.445 2.715 ;
        RECT 1.275 1.765 1.445 2.545 ;
        RECT 1.815 2.545 2.605 2.715 ;
        RECT 1.815 1.765 1.985 2.545 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 2.275 2.275 3.065 2.445 ;
        RECT 1.275 1.595 3.145 1.765 ;
        RECT 1.815 1.185 1.985 1.595 ;
        RECT 0.115 1.015 1.985 1.185 ;
  END
END AN2D1_3

#--------EOF---------

MACRO AO21D1
  CLASS CORE ;
  FOREIGN AO21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.105 0.905 2.445 ;
        RECT 0.655 1.935 0.985 2.105 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.105 3.065 2.445 ;
        RECT 2.815 1.935 3.145 2.105 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 4.435 2.545 4.765 2.715 ;
        RECT 4.515 1.185 4.685 2.545 ;
        RECT 4.435 1.015 4.765 1.185 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 0.000 -0.085 6.460 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.460 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 6.460 4.165 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 6.460 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 6.640 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 5.955 1.395 ;
      LAYER li1 ;
        RECT 0.115 2.885 2.605 3.055 ;
        RECT 0.195 2.545 1.525 2.715 ;
        RECT 0.195 1.765 0.365 2.545 ;
        RECT 0.195 1.595 4.225 1.765 ;
        RECT 0.195 1.185 0.365 1.595 ;
        RECT 3.435 1.185 3.605 1.595 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
  END
END AO21D1

#--------EOF---------

MACRO AO21D1_1
  CLASS CORE ;
  FOREIGN AO21D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.435 1.765 3.605 2.105 ;
        RECT 3.355 1.595 3.685 1.765 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 5.515 2.545 5.845 2.715 ;
        RECT 5.595 1.185 5.765 2.545 ;
        RECT 5.515 1.015 5.845 1.185 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 0.000 -0.085 6.460 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.460 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 6.460 4.165 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 6.460 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 6.640 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 5.955 1.395 ;
      LAYER li1 ;
        RECT 0.115 2.885 4.145 3.055 ;
        RECT 3.975 1.765 4.145 2.885 ;
        RECT 3.975 1.595 5.305 1.765 ;
        RECT 3.975 1.185 4.145 1.595 ;
        RECT 2.275 1.015 4.145 1.185 ;
        RECT 1.195 2.545 3.685 2.715 ;
  END
END AO21D1_1

#--------EOF---------

MACRO AO21D1_2
  CLASS CORE ;
  FOREIGN AO21D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.815 1.935 3.145 2.105 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 4.435 2.545 5.225 2.715 ;
        RECT 5.055 1.185 5.225 2.545 ;
        RECT 4.435 1.015 5.225 1.185 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 3.435 0.085 3.605 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 0.000 -0.085 6.460 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.460 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 6.460 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 6.460 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 6.640 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 5.955 1.395 ;
      LAYER li1 ;
        RECT 1.195 2.545 3.685 2.715 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 1.275 2.275 4.225 2.445 ;
        RECT 1.275 1.185 1.445 2.275 ;
        RECT 2.355 1.765 2.525 2.275 ;
        RECT 2.355 1.595 4.765 1.765 ;
        RECT 1.195 1.015 1.525 1.185 ;
  END
END AO21D1_2

#--------EOF---------

MACRO AO21D1_3
  CLASS CORE ;
  FOREIGN AO21D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 1.765 3.065 2.105 ;
        RECT 2.815 1.595 3.145 1.765 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 4.435 2.545 4.765 2.715 ;
        RECT 4.515 1.185 4.685 2.545 ;
        RECT 4.435 1.015 4.765 1.185 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 0.000 -0.085 6.460 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.460 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 6.460 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 6.460 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 6.640 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 5.955 1.395 ;
      LAYER li1 ;
        RECT 1.195 2.545 3.685 2.715 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 0.195 2.275 4.145 2.445 ;
        RECT 0.195 1.185 0.365 2.275 ;
        RECT 3.975 1.765 4.145 2.275 ;
        RECT 3.895 1.595 4.225 1.765 ;
        RECT 3.975 1.185 4.145 1.595 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 3.355 1.015 4.145 1.185 ;
  END
END AO21D1_3

#--------EOF---------

MACRO AOI21D1
  CLASS CORE ;
  FOREIGN AOI21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.080 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.074500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.545 2.605 2.715 ;
        RECT 1.275 1.765 1.445 2.545 ;
        RECT 1.275 1.595 2.525 1.765 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 2.275 1.015 2.605 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 1.765 3.065 2.105 ;
        RECT 2.815 1.595 3.145 1.765 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 3.435 0.085 3.605 1.015 ;
        RECT 0.000 -0.085 4.080 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.080 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 4.080 4.165 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 3.355 2.885 3.685 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 4.080 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 4.260 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 3.795 1.395 ;
  END
END AOI21D1

#--------EOF---------

MACRO AOI21D1_1
  CLASS CORE ;
  FOREIGN AOI21D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.080 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.074500 ;
    PORT
      LAYER li1 ;
        RECT 1.195 2.545 3.685 2.715 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 1.275 2.275 2.525 2.445 ;
        RECT 1.275 1.185 1.445 2.275 ;
        RECT 1.195 1.015 1.525 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 1.765 3.065 2.105 ;
        RECT 2.815 1.595 3.145 1.765 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 3.435 0.085 3.605 1.015 ;
        RECT 0.000 -0.085 4.080 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.080 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 4.080 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 4.080 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 4.260 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 3.795 1.395 ;
  END
END AOI21D1_1

#--------EOF---------

MACRO AOI21D1_2
  CLASS CORE ;
  FOREIGN AOI21D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.553000 ;
    PORT
      LAYER li1 ;
        RECT 1.275 3.605 3.605 3.775 ;
        RECT 1.275 3.055 1.445 3.605 ;
        RECT 3.435 3.055 3.605 3.605 ;
        RECT 0.115 2.885 3.065 3.055 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 2.895 2.715 3.065 2.885 ;
        RECT 2.275 2.545 3.065 2.715 ;
        RECT 2.895 1.185 3.065 2.545 ;
        RECT 2.275 1.015 3.685 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.975 1.765 4.145 2.105 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 0.000 -0.085 5.440 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 5.440 4.165 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 5.440 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 5.620 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 4.875 1.395 ;
  END
END AOI21D1_2

#--------EOF---------

MACRO AOI21D1_3
  CLASS CORE ;
  FOREIGN AOI21D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.553000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 1.195 2.545 3.685 2.715 ;
        RECT 0.195 2.445 0.365 2.545 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 0.195 2.275 2.525 2.445 ;
        RECT 0.195 1.185 0.365 2.275 ;
        RECT 2.355 1.765 2.525 2.275 ;
        RECT 2.355 1.595 3.605 1.765 ;
        RECT 3.435 1.185 3.605 1.595 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.975 1.765 4.145 2.105 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 0.000 -0.085 5.440 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 5.440 4.165 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 5.440 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 5.620 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 4.875 1.395 ;
  END
END AOI21D1_3

#--------EOF---------

MACRO BUFFD1
  CLASS CORE ;
  FOREIGN BUFFD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.060 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 0.195 1.185 0.365 2.545 ;
        RECT 0.115 1.015 0.445 1.185 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138000 ;
    PORT
      LAYER li1 ;
        RECT 1.735 2.545 2.065 2.715 ;
        RECT 1.815 1.765 1.985 2.545 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 0.000 -0.085 3.060 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.060 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 3.060 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 3.060 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 3.240 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 2.715 1.395 ;
        RECT 0.005 0.485 1.635 0.715 ;
      LAYER li1 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 2.355 2.445 2.525 2.885 ;
        RECT 2.275 2.275 2.605 2.445 ;
        RECT 2.275 1.595 2.605 1.765 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 2.275 1.015 2.605 1.185 ;
  END
END BUFFD1

#--------EOF---------

MACRO BUFFD1_1
  CLASS CORE ;
  FOREIGN BUFFD1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.060 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 2.275 2.545 2.605 2.715 ;
        RECT 2.355 1.185 2.525 2.545 ;
        RECT 2.275 1.015 2.605 1.185 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 0.000 -0.085 3.060 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.060 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 3.060 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 3.060 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 3.240 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 2.715 1.395 ;
        RECT 1.085 0.485 2.715 0.715 ;
      LAYER li1 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 0.195 1.185 0.365 2.885 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 0.195 0.475 0.365 1.015 ;
        RECT 0.115 0.305 0.445 0.475 ;
  END
END BUFFD1_1

#--------EOF---------

MACRO DFCNQD1
  CLASS CORE ;
  FOREIGN DFCNQD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.380 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.173250 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END d
  PIN cdn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.358500 ;
    PORT
      LAYER li1 ;
        RECT 5.055 2.105 5.225 2.445 ;
        RECT 4.975 1.935 5.305 2.105 ;
    END
  END cdn
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138000 ;
    PORT
      LAYER li1 ;
        RECT 18.015 1.765 18.185 2.105 ;
        RECT 17.935 1.595 18.265 1.765 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 16.315 2.545 16.645 2.715 ;
        RECT 16.395 1.185 16.565 2.545 ;
        RECT 16.315 1.015 16.645 1.185 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 10.915 1.015 11.245 1.185 ;
        RECT 15.235 1.015 15.565 1.185 ;
        RECT 18.475 1.015 18.805 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 10.995 0.085 11.165 1.015 ;
        RECT 15.315 0.085 15.485 1.015 ;
        RECT 18.555 0.085 18.725 1.015 ;
        RECT 0.000 -0.085 19.380 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
        RECT 10.965 -0.085 11.135 0.085 ;
        RECT 11.305 -0.085 11.475 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 11.985 -0.085 12.155 0.085 ;
        RECT 12.325 -0.085 12.495 0.085 ;
        RECT 12.665 -0.085 12.835 0.085 ;
        RECT 13.005 -0.085 13.175 0.085 ;
        RECT 13.345 -0.085 13.515 0.085 ;
        RECT 13.685 -0.085 13.855 0.085 ;
        RECT 14.025 -0.085 14.195 0.085 ;
        RECT 14.365 -0.085 14.535 0.085 ;
        RECT 14.705 -0.085 14.875 0.085 ;
        RECT 15.045 -0.085 15.215 0.085 ;
        RECT 15.385 -0.085 15.555 0.085 ;
        RECT 15.725 -0.085 15.895 0.085 ;
        RECT 16.065 -0.085 16.235 0.085 ;
        RECT 16.405 -0.085 16.575 0.085 ;
        RECT 16.745 -0.085 16.915 0.085 ;
        RECT 17.085 -0.085 17.255 0.085 ;
        RECT 17.425 -0.085 17.595 0.085 ;
        RECT 17.765 -0.085 17.935 0.085 ;
        RECT 18.105 -0.085 18.275 0.085 ;
        RECT 18.445 -0.085 18.615 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.125 -0.085 19.295 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 19.380 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 19.380 4.165 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 10.995 3.055 11.165 3.995 ;
        RECT 15.315 3.055 15.485 3.995 ;
        RECT 18.555 3.055 18.725 3.995 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
        RECT 10.915 2.885 11.245 3.055 ;
        RECT 15.235 2.885 15.565 3.055 ;
        RECT 18.475 2.885 18.805 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
        RECT 10.965 3.995 11.135 4.165 ;
        RECT 11.305 3.995 11.475 4.165 ;
        RECT 11.645 3.995 11.815 4.165 ;
        RECT 11.985 3.995 12.155 4.165 ;
        RECT 12.325 3.995 12.495 4.165 ;
        RECT 12.665 3.995 12.835 4.165 ;
        RECT 13.005 3.995 13.175 4.165 ;
        RECT 13.345 3.995 13.515 4.165 ;
        RECT 13.685 3.995 13.855 4.165 ;
        RECT 14.025 3.995 14.195 4.165 ;
        RECT 14.365 3.995 14.535 4.165 ;
        RECT 14.705 3.995 14.875 4.165 ;
        RECT 15.045 3.995 15.215 4.165 ;
        RECT 15.385 3.995 15.555 4.165 ;
        RECT 15.725 3.995 15.895 4.165 ;
        RECT 16.065 3.995 16.235 4.165 ;
        RECT 16.405 3.995 16.575 4.165 ;
        RECT 16.745 3.995 16.915 4.165 ;
        RECT 17.085 3.995 17.255 4.165 ;
        RECT 17.425 3.995 17.595 4.165 ;
        RECT 17.765 3.995 17.935 4.165 ;
        RECT 18.105 3.995 18.275 4.165 ;
        RECT 18.445 3.995 18.615 4.165 ;
        RECT 18.785 3.995 18.955 4.165 ;
        RECT 19.125 3.995 19.295 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 19.380 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 19.560 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 18.915 1.395 ;
        RECT 5.405 0.680 10.275 0.715 ;
        RECT 5.405 0.485 8.115 0.680 ;
        RECT 15.125 0.485 16.755 0.715 ;
      LAYER li1 ;
        RECT 9.835 3.605 10.165 3.775 ;
        RECT 9.915 3.055 10.085 3.605 ;
        RECT 9.835 2.885 10.165 3.055 ;
        RECT 14.695 2.275 15.025 2.445 ;
        RECT 9.835 1.015 10.165 1.185 ;
        RECT 9.915 0.475 10.085 1.015 ;
        RECT 14.775 0.475 14.945 2.275 ;
        RECT 9.835 0.305 10.165 0.475 ;
        RECT 14.695 0.305 15.025 0.475 ;
        RECT 14.155 2.885 14.485 3.055 ;
        RECT 9.835 1.935 11.785 2.105 ;
        RECT 14.235 1.185 14.405 2.885 ;
        RECT 13.615 1.015 14.485 1.185 ;
        RECT 13.075 2.885 13.405 3.055 ;
        RECT 8.755 2.545 9.085 2.715 ;
        RECT 8.835 2.445 9.005 2.545 ;
        RECT 8.755 2.275 12.245 2.445 ;
        RECT 12.075 1.765 12.245 2.275 ;
        RECT 13.155 1.765 13.325 2.885 ;
        RECT 12.075 1.595 13.325 1.765 ;
        RECT 13.155 1.185 13.325 1.595 ;
        RECT 8.215 1.015 9.085 1.185 ;
        RECT 13.075 1.015 13.405 1.185 ;
        RECT 0.115 2.885 3.065 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
        RECT 1.275 1.765 1.445 2.885 ;
        RECT 2.895 2.715 3.065 2.885 ;
        RECT 4.515 2.715 4.685 2.885 ;
        RECT 2.895 2.545 4.685 2.715 ;
        RECT 1.275 1.595 10.705 1.765 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 2.275 1.015 2.605 1.185 ;
  END
END DFCNQD1

#--------EOF---------

MACRO DFCNQD1_1
  CLASS CORE ;
  FOREIGN DFCNQD1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.380 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.173250 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END d
  PIN cdn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.358500 ;
    PORT
      LAYER li1 ;
        RECT 5.055 2.105 5.225 2.445 ;
        RECT 4.975 1.935 5.305 2.105 ;
    END
  END cdn
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138000 ;
    PORT
      LAYER li1 ;
        RECT 18.015 1.765 18.185 2.105 ;
        RECT 17.935 1.595 18.265 1.765 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 14.155 2.545 14.485 2.715 ;
        RECT 14.235 1.185 14.405 2.545 ;
        RECT 14.155 1.015 14.485 1.185 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 10.915 1.015 11.245 1.185 ;
        RECT 15.235 1.015 15.565 1.185 ;
        RECT 18.475 1.015 18.805 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 10.995 0.085 11.165 1.015 ;
        RECT 15.315 0.085 15.485 1.015 ;
        RECT 18.555 0.085 18.725 1.015 ;
        RECT 0.000 -0.085 19.380 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
        RECT 10.965 -0.085 11.135 0.085 ;
        RECT 11.305 -0.085 11.475 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 11.985 -0.085 12.155 0.085 ;
        RECT 12.325 -0.085 12.495 0.085 ;
        RECT 12.665 -0.085 12.835 0.085 ;
        RECT 13.005 -0.085 13.175 0.085 ;
        RECT 13.345 -0.085 13.515 0.085 ;
        RECT 13.685 -0.085 13.855 0.085 ;
        RECT 14.025 -0.085 14.195 0.085 ;
        RECT 14.365 -0.085 14.535 0.085 ;
        RECT 14.705 -0.085 14.875 0.085 ;
        RECT 15.045 -0.085 15.215 0.085 ;
        RECT 15.385 -0.085 15.555 0.085 ;
        RECT 15.725 -0.085 15.895 0.085 ;
        RECT 16.065 -0.085 16.235 0.085 ;
        RECT 16.405 -0.085 16.575 0.085 ;
        RECT 16.745 -0.085 16.915 0.085 ;
        RECT 17.085 -0.085 17.255 0.085 ;
        RECT 17.425 -0.085 17.595 0.085 ;
        RECT 17.765 -0.085 17.935 0.085 ;
        RECT 18.105 -0.085 18.275 0.085 ;
        RECT 18.445 -0.085 18.615 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.125 -0.085 19.295 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 19.380 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 19.380 4.165 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 10.995 3.055 11.165 3.995 ;
        RECT 15.315 3.055 15.485 3.995 ;
        RECT 18.555 3.055 18.725 3.995 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
        RECT 10.915 2.885 11.245 3.055 ;
        RECT 15.235 2.885 15.565 3.055 ;
        RECT 18.475 2.885 18.805 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
        RECT 10.965 3.995 11.135 4.165 ;
        RECT 11.305 3.995 11.475 4.165 ;
        RECT 11.645 3.995 11.815 4.165 ;
        RECT 11.985 3.995 12.155 4.165 ;
        RECT 12.325 3.995 12.495 4.165 ;
        RECT 12.665 3.995 12.835 4.165 ;
        RECT 13.005 3.995 13.175 4.165 ;
        RECT 13.345 3.995 13.515 4.165 ;
        RECT 13.685 3.995 13.855 4.165 ;
        RECT 14.025 3.995 14.195 4.165 ;
        RECT 14.365 3.995 14.535 4.165 ;
        RECT 14.705 3.995 14.875 4.165 ;
        RECT 15.045 3.995 15.215 4.165 ;
        RECT 15.385 3.995 15.555 4.165 ;
        RECT 15.725 3.995 15.895 4.165 ;
        RECT 16.065 3.995 16.235 4.165 ;
        RECT 16.405 3.995 16.575 4.165 ;
        RECT 16.745 3.995 16.915 4.165 ;
        RECT 17.085 3.995 17.255 4.165 ;
        RECT 17.425 3.995 17.595 4.165 ;
        RECT 17.765 3.995 17.935 4.165 ;
        RECT 18.105 3.995 18.275 4.165 ;
        RECT 18.445 3.995 18.615 4.165 ;
        RECT 18.785 3.995 18.955 4.165 ;
        RECT 19.125 3.995 19.295 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 19.380 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 19.560 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 18.915 1.395 ;
        RECT 5.405 0.680 10.275 0.715 ;
        RECT 5.405 0.485 8.115 0.680 ;
        RECT 14.045 0.485 15.675 0.715 ;
      LAYER li1 ;
        RECT 9.835 3.605 10.165 3.775 ;
        RECT 9.915 3.055 10.085 3.605 ;
        RECT 9.835 2.885 10.165 3.055 ;
        RECT 13.615 2.275 13.945 2.445 ;
        RECT 9.835 1.015 10.165 1.185 ;
        RECT 9.915 0.475 10.085 1.015 ;
        RECT 13.695 0.475 13.865 2.275 ;
        RECT 9.835 0.305 10.165 0.475 ;
        RECT 11.455 0.305 13.865 0.475 ;
        RECT 16.315 2.885 16.645 3.055 ;
        RECT 9.835 1.935 11.785 2.105 ;
        RECT 16.395 1.765 16.565 2.885 ;
        RECT 16.315 1.595 16.645 1.765 ;
        RECT 16.395 1.185 16.565 1.595 ;
        RECT 16.315 1.015 16.645 1.185 ;
        RECT 13.075 2.885 13.405 3.055 ;
        RECT 8.755 2.545 9.085 2.715 ;
        RECT 8.835 2.445 9.005 2.545 ;
        RECT 8.755 2.275 12.245 2.445 ;
        RECT 12.075 1.765 12.245 2.275 ;
        RECT 13.155 1.765 13.325 2.885 ;
        RECT 12.075 1.595 13.325 1.765 ;
        RECT 13.155 1.185 13.325 1.595 ;
        RECT 8.215 1.015 9.085 1.185 ;
        RECT 13.075 1.015 13.405 1.185 ;
        RECT 0.115 2.885 3.065 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
        RECT 1.275 1.765 1.445 2.885 ;
        RECT 2.895 2.715 3.065 2.885 ;
        RECT 4.515 2.715 4.685 2.885 ;
        RECT 2.895 2.545 4.685 2.715 ;
        RECT 1.275 1.595 10.705 1.765 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 2.275 1.015 2.605 1.185 ;
  END
END DFCNQD1_1

#--------EOF---------

MACRO DFCNQD1_2
  CLASS CORE ;
  FOREIGN DFCNQD1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.380 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.173250 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END d
  PIN cdn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.358500 ;
    PORT
      LAYER li1 ;
        RECT 5.055 2.715 5.225 3.055 ;
        RECT 4.975 2.545 5.305 2.715 ;
    END
  END cdn
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138000 ;
    PORT
      LAYER li1 ;
        RECT 18.015 1.765 18.185 2.105 ;
        RECT 17.935 1.595 18.265 1.765 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 16.315 2.545 16.645 2.715 ;
        RECT 16.395 1.185 16.565 2.545 ;
        RECT 16.315 1.015 16.645 1.185 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 9.835 1.015 10.165 1.185 ;
        RECT 15.235 1.015 15.565 1.185 ;
        RECT 18.475 1.015 18.805 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 9.915 0.085 10.085 1.015 ;
        RECT 15.315 0.085 15.485 1.015 ;
        RECT 18.555 0.085 18.725 1.015 ;
        RECT 0.000 -0.085 19.380 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
        RECT 10.965 -0.085 11.135 0.085 ;
        RECT 11.305 -0.085 11.475 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 11.985 -0.085 12.155 0.085 ;
        RECT 12.325 -0.085 12.495 0.085 ;
        RECT 12.665 -0.085 12.835 0.085 ;
        RECT 13.005 -0.085 13.175 0.085 ;
        RECT 13.345 -0.085 13.515 0.085 ;
        RECT 13.685 -0.085 13.855 0.085 ;
        RECT 14.025 -0.085 14.195 0.085 ;
        RECT 14.365 -0.085 14.535 0.085 ;
        RECT 14.705 -0.085 14.875 0.085 ;
        RECT 15.045 -0.085 15.215 0.085 ;
        RECT 15.385 -0.085 15.555 0.085 ;
        RECT 15.725 -0.085 15.895 0.085 ;
        RECT 16.065 -0.085 16.235 0.085 ;
        RECT 16.405 -0.085 16.575 0.085 ;
        RECT 16.745 -0.085 16.915 0.085 ;
        RECT 17.085 -0.085 17.255 0.085 ;
        RECT 17.425 -0.085 17.595 0.085 ;
        RECT 17.765 -0.085 17.935 0.085 ;
        RECT 18.105 -0.085 18.275 0.085 ;
        RECT 18.445 -0.085 18.615 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.125 -0.085 19.295 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 19.380 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 19.380 4.165 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 9.915 3.055 10.085 3.995 ;
        RECT 15.315 3.055 15.485 3.995 ;
        RECT 18.555 3.055 18.725 3.995 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
        RECT 9.835 2.885 10.165 3.055 ;
        RECT 15.235 2.885 15.565 3.055 ;
        RECT 18.475 2.885 18.805 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
        RECT 10.965 3.995 11.135 4.165 ;
        RECT 11.305 3.995 11.475 4.165 ;
        RECT 11.645 3.995 11.815 4.165 ;
        RECT 11.985 3.995 12.155 4.165 ;
        RECT 12.325 3.995 12.495 4.165 ;
        RECT 12.665 3.995 12.835 4.165 ;
        RECT 13.005 3.995 13.175 4.165 ;
        RECT 13.345 3.995 13.515 4.165 ;
        RECT 13.685 3.995 13.855 4.165 ;
        RECT 14.025 3.995 14.195 4.165 ;
        RECT 14.365 3.995 14.535 4.165 ;
        RECT 14.705 3.995 14.875 4.165 ;
        RECT 15.045 3.995 15.215 4.165 ;
        RECT 15.385 3.995 15.555 4.165 ;
        RECT 15.725 3.995 15.895 4.165 ;
        RECT 16.065 3.995 16.235 4.165 ;
        RECT 16.405 3.995 16.575 4.165 ;
        RECT 16.745 3.995 16.915 4.165 ;
        RECT 17.085 3.995 17.255 4.165 ;
        RECT 17.425 3.995 17.595 4.165 ;
        RECT 17.765 3.995 17.935 4.165 ;
        RECT 18.105 3.995 18.275 4.165 ;
        RECT 18.445 3.995 18.615 4.165 ;
        RECT 18.785 3.995 18.955 4.165 ;
        RECT 19.125 3.995 19.295 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 19.380 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 19.560 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 18.915 1.395 ;
        RECT 5.405 0.485 8.115 0.715 ;
        RECT 11.885 0.680 13.515 0.715 ;
        RECT 15.125 0.485 16.755 0.715 ;
      LAYER li1 ;
        RECT 12.535 3.605 12.865 3.775 ;
        RECT 8.215 2.885 9.085 3.055 ;
        RECT 12.615 2.715 12.785 3.605 ;
        RECT 12.615 2.545 13.405 2.715 ;
        RECT 3.895 1.935 8.005 2.105 ;
        RECT 12.615 1.185 12.785 2.545 ;
        RECT 8.215 1.015 9.085 1.185 ;
        RECT 12.615 1.015 13.405 1.185 ;
        RECT 14.155 2.885 14.485 3.055 ;
        RECT 11.455 2.545 11.785 2.715 ;
        RECT 11.535 2.445 11.705 2.545 ;
        RECT 4.435 2.275 11.705 2.445 ;
        RECT 14.235 1.765 14.405 2.885 ;
        RECT 14.155 1.595 14.485 1.765 ;
        RECT 14.235 1.185 14.405 1.595 ;
        RECT 14.155 1.015 14.485 1.185 ;
        RECT 11.995 2.885 12.325 3.055 ;
        RECT 12.075 1.185 12.245 2.885 ;
        RECT 11.995 1.015 12.325 1.185 ;
        RECT 12.075 0.475 12.245 1.015 ;
        RECT 11.995 0.305 12.325 0.475 ;
        RECT 0.115 2.885 3.065 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
        RECT 1.275 1.765 1.445 2.885 ;
        RECT 2.895 2.715 3.065 2.885 ;
        RECT 4.515 2.715 4.685 2.885 ;
        RECT 2.895 2.545 4.685 2.715 ;
        RECT 1.275 1.595 9.625 1.765 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 2.275 1.015 2.605 1.185 ;
  END
END DFCNQD1_2

#--------EOF---------

MACRO DFCNQD1_3
  CLASS CORE ;
  FOREIGN DFCNQD1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.380 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.173250 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END d
  PIN cdn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.358500 ;
    PORT
      LAYER li1 ;
        RECT 5.055 2.715 5.225 3.055 ;
        RECT 4.975 2.545 5.305 2.715 ;
    END
  END cdn
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138000 ;
    PORT
      LAYER li1 ;
        RECT 18.015 1.765 18.185 2.105 ;
        RECT 17.935 1.595 18.265 1.765 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 14.155 2.545 14.485 2.715 ;
        RECT 14.235 1.185 14.405 2.545 ;
        RECT 14.155 1.015 14.485 1.185 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 9.835 1.015 10.165 1.185 ;
        RECT 15.235 1.015 15.565 1.185 ;
        RECT 18.475 1.015 18.805 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 9.915 0.085 10.085 1.015 ;
        RECT 15.315 0.085 15.485 1.015 ;
        RECT 18.555 0.085 18.725 1.015 ;
        RECT 0.000 -0.085 19.380 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
        RECT 10.965 -0.085 11.135 0.085 ;
        RECT 11.305 -0.085 11.475 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 11.985 -0.085 12.155 0.085 ;
        RECT 12.325 -0.085 12.495 0.085 ;
        RECT 12.665 -0.085 12.835 0.085 ;
        RECT 13.005 -0.085 13.175 0.085 ;
        RECT 13.345 -0.085 13.515 0.085 ;
        RECT 13.685 -0.085 13.855 0.085 ;
        RECT 14.025 -0.085 14.195 0.085 ;
        RECT 14.365 -0.085 14.535 0.085 ;
        RECT 14.705 -0.085 14.875 0.085 ;
        RECT 15.045 -0.085 15.215 0.085 ;
        RECT 15.385 -0.085 15.555 0.085 ;
        RECT 15.725 -0.085 15.895 0.085 ;
        RECT 16.065 -0.085 16.235 0.085 ;
        RECT 16.405 -0.085 16.575 0.085 ;
        RECT 16.745 -0.085 16.915 0.085 ;
        RECT 17.085 -0.085 17.255 0.085 ;
        RECT 17.425 -0.085 17.595 0.085 ;
        RECT 17.765 -0.085 17.935 0.085 ;
        RECT 18.105 -0.085 18.275 0.085 ;
        RECT 18.445 -0.085 18.615 0.085 ;
        RECT 18.785 -0.085 18.955 0.085 ;
        RECT 19.125 -0.085 19.295 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 19.380 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 19.380 4.165 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 9.915 3.055 10.085 3.995 ;
        RECT 15.315 3.055 15.485 3.995 ;
        RECT 18.555 3.055 18.725 3.995 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
        RECT 9.835 2.885 10.165 3.055 ;
        RECT 15.235 2.885 15.565 3.055 ;
        RECT 18.475 2.885 18.805 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
        RECT 10.965 3.995 11.135 4.165 ;
        RECT 11.305 3.995 11.475 4.165 ;
        RECT 11.645 3.995 11.815 4.165 ;
        RECT 11.985 3.995 12.155 4.165 ;
        RECT 12.325 3.995 12.495 4.165 ;
        RECT 12.665 3.995 12.835 4.165 ;
        RECT 13.005 3.995 13.175 4.165 ;
        RECT 13.345 3.995 13.515 4.165 ;
        RECT 13.685 3.995 13.855 4.165 ;
        RECT 14.025 3.995 14.195 4.165 ;
        RECT 14.365 3.995 14.535 4.165 ;
        RECT 14.705 3.995 14.875 4.165 ;
        RECT 15.045 3.995 15.215 4.165 ;
        RECT 15.385 3.995 15.555 4.165 ;
        RECT 15.725 3.995 15.895 4.165 ;
        RECT 16.065 3.995 16.235 4.165 ;
        RECT 16.405 3.995 16.575 4.165 ;
        RECT 16.745 3.995 16.915 4.165 ;
        RECT 17.085 3.995 17.255 4.165 ;
        RECT 17.425 3.995 17.595 4.165 ;
        RECT 17.765 3.995 17.935 4.165 ;
        RECT 18.105 3.995 18.275 4.165 ;
        RECT 18.445 3.995 18.615 4.165 ;
        RECT 18.785 3.995 18.955 4.165 ;
        RECT 19.125 3.995 19.295 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 19.380 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 19.560 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 18.915 1.395 ;
        RECT 5.405 0.485 8.115 0.715 ;
        RECT 11.885 0.680 15.675 0.715 ;
        RECT 14.045 0.485 15.675 0.680 ;
      LAYER li1 ;
        RECT 12.535 3.605 12.865 3.775 ;
        RECT 8.215 2.885 9.085 3.055 ;
        RECT 12.615 2.715 12.785 3.605 ;
        RECT 12.615 2.545 13.405 2.715 ;
        RECT 3.895 1.935 8.005 2.105 ;
        RECT 12.615 1.185 12.785 2.545 ;
        RECT 8.215 1.015 9.085 1.185 ;
        RECT 12.615 1.015 13.405 1.185 ;
        RECT 16.315 2.885 16.645 3.055 ;
        RECT 11.455 2.545 11.785 2.715 ;
        RECT 11.535 2.445 11.705 2.545 ;
        RECT 4.435 2.275 11.705 2.445 ;
        RECT 16.395 1.765 16.565 2.885 ;
        RECT 16.315 1.595 16.645 1.765 ;
        RECT 16.395 1.185 16.565 1.595 ;
        RECT 16.315 1.015 16.645 1.185 ;
        RECT 11.995 2.885 12.325 3.055 ;
        RECT 12.075 1.185 12.245 2.885 ;
        RECT 11.995 1.015 12.325 1.185 ;
        RECT 12.075 0.475 12.245 1.015 ;
        RECT 11.995 0.305 12.325 0.475 ;
        RECT 0.115 2.885 3.065 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
        RECT 1.275 1.765 1.445 2.885 ;
        RECT 2.895 2.715 3.065 2.885 ;
        RECT 4.515 2.715 4.685 2.885 ;
        RECT 2.895 2.545 4.685 2.715 ;
        RECT 1.275 1.595 9.625 1.765 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 2.275 1.015 2.605 1.185 ;
  END
END DFCNQD1_3

#--------EOF---------

MACRO DFQD1
  CLASS CORE ;
  FOREIGN DFQD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.980 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156750 ;
    PORT
      LAYER li1 ;
        RECT 2.815 2.545 3.145 2.715 ;
        RECT 2.895 1.765 3.065 2.545 ;
        RECT 2.815 1.595 3.145 1.765 ;
    END
  END d
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 14.155 2.545 14.485 2.715 ;
        RECT 14.235 1.185 14.405 2.545 ;
        RECT 14.155 1.015 14.485 1.185 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 11.995 1.015 12.325 1.185 ;
        RECT 15.235 1.015 15.565 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 12.075 0.085 12.245 1.015 ;
        RECT 15.315 0.085 15.485 1.015 ;
        RECT 0.000 -0.085 15.980 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
        RECT 10.965 -0.085 11.135 0.085 ;
        RECT 11.305 -0.085 11.475 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 11.985 -0.085 12.155 0.085 ;
        RECT 12.325 -0.085 12.495 0.085 ;
        RECT 12.665 -0.085 12.835 0.085 ;
        RECT 13.005 -0.085 13.175 0.085 ;
        RECT 13.345 -0.085 13.515 0.085 ;
        RECT 13.685 -0.085 13.855 0.085 ;
        RECT 14.025 -0.085 14.195 0.085 ;
        RECT 14.365 -0.085 14.535 0.085 ;
        RECT 14.705 -0.085 14.875 0.085 ;
        RECT 15.045 -0.085 15.215 0.085 ;
        RECT 15.385 -0.085 15.555 0.085 ;
        RECT 15.725 -0.085 15.895 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 15.980 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 15.980 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 12.075 3.055 12.245 3.995 ;
        RECT 15.315 3.055 15.485 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
        RECT 11.995 2.885 12.325 3.055 ;
        RECT 15.235 2.885 15.565 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
        RECT 10.965 3.995 11.135 4.165 ;
        RECT 11.305 3.995 11.475 4.165 ;
        RECT 11.645 3.995 11.815 4.165 ;
        RECT 11.985 3.995 12.155 4.165 ;
        RECT 12.325 3.995 12.495 4.165 ;
        RECT 12.665 3.995 12.835 4.165 ;
        RECT 13.005 3.995 13.175 4.165 ;
        RECT 13.345 3.995 13.515 4.165 ;
        RECT 13.685 3.995 13.855 4.165 ;
        RECT 14.025 3.995 14.195 4.165 ;
        RECT 14.365 3.995 14.535 4.165 ;
        RECT 14.705 3.995 14.875 4.165 ;
        RECT 15.045 3.995 15.215 4.165 ;
        RECT 15.385 3.995 15.555 4.165 ;
        RECT 15.725 3.995 15.895 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 15.980 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 16.160 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 15.675 1.395 ;
        RECT 0.005 0.485 1.635 0.715 ;
        RECT 5.405 0.710 9.195 0.715 ;
        RECT 5.405 0.485 7.035 0.710 ;
        RECT 11.885 0.485 15.675 0.715 ;
      LAYER li1 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 0.195 1.185 0.365 2.545 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 0.195 0.475 0.365 1.015 ;
        RECT 0.115 0.305 0.445 0.475 ;
        RECT 9.835 2.545 10.165 2.715 ;
        RECT 9.915 2.445 10.085 2.545 ;
        RECT 9.915 2.275 12.865 2.445 ;
        RECT 9.915 1.185 10.085 2.275 ;
        RECT 9.835 1.015 10.165 1.185 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 3.435 2.105 3.605 2.885 ;
        RECT 3.435 1.935 8.545 2.105 ;
        RECT 3.435 1.185 3.605 1.935 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 1.735 3.605 4.225 3.775 ;
        RECT 9.295 3.605 9.625 3.775 ;
        RECT 3.975 2.715 4.145 3.605 ;
        RECT 3.975 2.545 7.465 2.715 ;
        RECT 3.975 2.445 4.145 2.545 ;
        RECT 3.895 2.275 4.225 2.445 ;
        RECT 9.375 1.765 9.545 3.605 ;
        RECT 9.295 1.595 9.625 1.765 ;
        RECT 6.595 1.015 7.465 1.185 ;
        RECT 8.755 2.885 9.085 3.055 ;
        RECT 8.835 1.765 9.005 2.885 ;
        RECT 4.975 1.595 9.005 1.765 ;
        RECT 8.835 1.185 9.005 1.595 ;
        RECT 8.755 1.015 9.085 1.185 ;
        RECT 11.455 2.545 13.405 2.715 ;
        RECT 13.155 1.765 13.325 2.545 ;
        RECT 13.075 1.595 13.405 1.765 ;
        RECT 13.155 1.185 13.325 1.595 ;
        RECT 13.075 1.015 13.405 1.185 ;
  END
END DFQD1

#--------EOF---------

MACRO DFQD1_1
  CLASS CORE ;
  FOREIGN DFQD1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.960 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156750 ;
    PORT
      LAYER li1 ;
        RECT 2.815 1.595 3.145 1.765 ;
        RECT 2.895 1.015 3.065 1.595 ;
    END
  END d
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.105 0.905 2.445 ;
        RECT 0.655 1.935 0.985 2.105 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 14.155 2.545 14.485 2.715 ;
        RECT 14.235 1.185 14.405 2.545 ;
        RECT 14.155 1.015 14.485 1.185 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 9.835 1.015 10.165 1.185 ;
        RECT 13.075 1.015 13.405 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 9.915 0.085 10.085 1.015 ;
        RECT 13.155 0.085 13.325 1.015 ;
        RECT 0.000 -0.085 14.960 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
        RECT 10.965 -0.085 11.135 0.085 ;
        RECT 11.305 -0.085 11.475 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 11.985 -0.085 12.155 0.085 ;
        RECT 12.325 -0.085 12.495 0.085 ;
        RECT 12.665 -0.085 12.835 0.085 ;
        RECT 13.005 -0.085 13.175 0.085 ;
        RECT 13.345 -0.085 13.515 0.085 ;
        RECT 13.685 -0.085 13.855 0.085 ;
        RECT 14.025 -0.085 14.195 0.085 ;
        RECT 14.365 -0.085 14.535 0.085 ;
        RECT 14.705 -0.085 14.875 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 14.960 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 14.960 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 9.915 3.055 10.085 3.995 ;
        RECT 13.155 3.055 13.325 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 9.835 2.885 10.165 3.055 ;
        RECT 13.075 2.885 13.405 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
        RECT 10.965 3.995 11.135 4.165 ;
        RECT 11.305 3.995 11.475 4.165 ;
        RECT 11.645 3.995 11.815 4.165 ;
        RECT 11.985 3.995 12.155 4.165 ;
        RECT 12.325 3.995 12.495 4.165 ;
        RECT 12.665 3.995 12.835 4.165 ;
        RECT 13.005 3.995 13.175 4.165 ;
        RECT 13.345 3.995 13.515 4.165 ;
        RECT 13.685 3.995 13.855 4.165 ;
        RECT 14.025 3.995 14.195 4.165 ;
        RECT 14.365 3.995 14.535 4.165 ;
        RECT 14.705 3.995 14.875 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 14.960 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 15.140 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 14.595 1.395 ;
        RECT 0.005 0.485 1.635 0.715 ;
        RECT 5.405 0.710 7.035 0.715 ;
        RECT 9.725 0.485 14.595 0.715 ;
      LAYER li1 ;
        RECT 0.115 3.605 0.445 3.775 ;
        RECT 8.755 3.605 9.085 3.775 ;
        RECT 0.195 2.715 0.365 3.605 ;
        RECT 7.215 2.885 8.465 3.055 ;
        RECT 0.115 2.545 4.225 2.715 ;
        RECT 0.195 1.765 0.365 2.545 ;
        RECT 7.215 2.105 7.385 2.885 ;
        RECT 8.295 2.715 8.465 2.885 ;
        RECT 8.215 2.545 8.545 2.715 ;
        RECT 8.835 2.445 9.005 3.605 ;
        RECT 11.995 2.545 12.325 2.715 ;
        RECT 8.215 2.275 9.005 2.445 ;
        RECT 12.075 2.105 12.245 2.545 ;
        RECT 1.735 1.935 12.245 2.105 ;
        RECT 7.215 1.765 7.385 1.935 ;
        RECT 0.195 1.595 2.065 1.765 ;
        RECT 7.135 1.595 7.465 1.765 ;
        RECT 0.195 1.185 0.365 1.595 ;
        RECT 12.075 1.185 12.245 1.935 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 11.995 1.015 12.325 1.185 ;
        RECT 7.675 2.545 8.005 2.715 ;
        RECT 7.755 2.445 7.925 2.545 ;
        RECT 7.675 2.275 8.005 2.445 ;
        RECT 7.675 1.595 10.705 1.765 ;
        RECT 7.755 1.185 7.925 1.595 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 3.355 2.885 5.225 3.055 ;
        RECT 5.055 2.715 5.225 2.885 ;
        RECT 5.055 2.545 6.385 2.715 ;
        RECT 3.435 1.595 6.385 1.765 ;
        RECT 3.435 1.185 3.605 1.595 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 6.595 2.885 6.925 3.055 ;
        RECT 6.675 2.445 6.845 2.885 ;
        RECT 4.975 2.275 6.925 2.445 ;
        RECT 6.595 1.595 6.925 1.765 ;
        RECT 6.675 1.185 6.845 1.595 ;
        RECT 6.595 1.015 6.925 1.185 ;
        RECT 9.295 2.545 11.245 2.715 ;
        RECT 10.915 1.015 11.245 1.185 ;
        RECT 10.995 0.475 11.165 1.015 ;
        RECT 10.915 0.305 11.245 0.475 ;
  END
END DFQD1_1

#--------EOF---------

MACRO DFQD1_2
  CLASS CORE ;
  FOREIGN DFQD1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.980 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156750 ;
    PORT
      LAYER li1 ;
        RECT 4.975 1.595 5.305 1.765 ;
        RECT 5.055 1.015 5.225 1.595 ;
    END
  END d
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.256500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 2.275 0.985 2.445 ;
        RECT 0.735 1.765 0.905 2.275 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 14.155 2.545 14.485 2.715 ;
        RECT 14.235 1.185 14.405 2.545 ;
        RECT 14.155 1.015 14.485 1.185 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 11.995 1.015 12.325 1.185 ;
        RECT 15.235 1.015 15.565 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 3.435 0.085 3.605 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 12.075 0.085 12.245 1.015 ;
        RECT 15.315 0.085 15.485 1.015 ;
        RECT 0.000 -0.085 15.980 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
        RECT 10.965 -0.085 11.135 0.085 ;
        RECT 11.305 -0.085 11.475 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 11.985 -0.085 12.155 0.085 ;
        RECT 12.325 -0.085 12.495 0.085 ;
        RECT 12.665 -0.085 12.835 0.085 ;
        RECT 13.005 -0.085 13.175 0.085 ;
        RECT 13.345 -0.085 13.515 0.085 ;
        RECT 13.685 -0.085 13.855 0.085 ;
        RECT 14.025 -0.085 14.195 0.085 ;
        RECT 14.365 -0.085 14.535 0.085 ;
        RECT 14.705 -0.085 14.875 0.085 ;
        RECT 15.045 -0.085 15.215 0.085 ;
        RECT 15.385 -0.085 15.555 0.085 ;
        RECT 15.725 -0.085 15.895 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 15.980 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 15.980 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 12.075 3.055 12.245 3.995 ;
        RECT 15.315 3.055 15.485 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
        RECT 11.995 2.885 12.325 3.055 ;
        RECT 15.235 2.885 15.565 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
        RECT 10.965 3.995 11.135 4.165 ;
        RECT 11.305 3.995 11.475 4.165 ;
        RECT 11.645 3.995 11.815 4.165 ;
        RECT 11.985 3.995 12.155 4.165 ;
        RECT 12.325 3.995 12.495 4.165 ;
        RECT 12.665 3.995 12.835 4.165 ;
        RECT 13.005 3.995 13.175 4.165 ;
        RECT 13.345 3.995 13.515 4.165 ;
        RECT 13.685 3.995 13.855 4.165 ;
        RECT 14.025 3.995 14.195 4.165 ;
        RECT 14.365 3.995 14.535 4.165 ;
        RECT 14.705 3.995 14.875 4.165 ;
        RECT 15.045 3.995 15.215 4.165 ;
        RECT 15.385 3.995 15.555 4.165 ;
        RECT 15.725 3.995 15.895 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 15.980 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 16.160 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 15.675 1.395 ;
        RECT 0.005 0.485 2.715 0.715 ;
        RECT 7.565 0.710 9.195 0.715 ;
        RECT 11.885 0.485 15.675 0.715 ;
      LAYER li1 ;
        RECT 0.115 2.545 6.385 2.715 ;
        RECT 0.115 1.935 0.445 2.105 ;
        RECT 0.195 1.185 0.365 1.935 ;
        RECT 1.815 1.765 1.985 2.545 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 2.355 2.275 6.385 2.445 ;
        RECT 9.295 2.275 9.625 2.445 ;
        RECT 10.375 2.275 10.705 2.445 ;
        RECT 1.735 1.595 2.065 1.765 ;
        RECT 2.355 1.185 2.525 2.275 ;
        RECT 9.375 2.105 9.545 2.275 ;
        RECT 3.895 1.935 9.545 2.105 ;
        RECT 10.455 1.765 10.625 2.275 ;
        RECT 10.375 1.595 10.705 1.765 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 9.835 2.545 12.785 2.715 ;
        RECT 9.915 1.185 10.085 2.545 ;
        RECT 12.615 2.445 12.785 2.545 ;
        RECT 12.535 2.275 12.865 2.445 ;
        RECT 9.835 1.015 10.165 1.185 ;
        RECT 5.515 3.605 5.845 3.775 ;
        RECT 5.595 3.055 5.765 3.605 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 5.595 1.595 8.545 1.765 ;
        RECT 5.595 1.185 5.765 1.595 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 8.755 2.885 9.085 3.055 ;
        RECT 8.835 2.715 9.005 2.885 ;
        RECT 7.135 2.545 9.005 2.715 ;
        RECT 8.835 2.445 9.005 2.545 ;
        RECT 8.755 2.275 9.085 2.445 ;
        RECT 8.755 1.595 9.085 1.765 ;
        RECT 8.835 1.185 9.005 1.595 ;
        RECT 8.755 1.015 9.085 1.185 ;
        RECT 13.075 3.605 13.405 3.775 ;
        RECT 13.155 3.055 13.325 3.605 ;
        RECT 13.075 2.885 13.405 3.055 ;
        RECT 13.075 2.545 13.405 2.715 ;
        RECT 13.155 1.185 13.325 2.545 ;
        RECT 13.075 1.015 13.405 1.185 ;
        RECT 13.155 0.475 13.325 1.015 ;
        RECT 13.075 0.305 13.405 0.475 ;
  END
END DFQD1_2

#--------EOF---------

MACRO DFQD1_3
  CLASS CORE ;
  FOREIGN DFQD1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.980 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156750 ;
    PORT
      LAYER li1 ;
        RECT 4.975 1.595 5.305 1.765 ;
        RECT 5.055 1.015 5.225 1.595 ;
    END
  END d
  PIN cp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END cp
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 14.155 2.545 14.485 2.715 ;
        RECT 14.235 1.185 14.405 2.545 ;
        RECT 14.155 1.015 14.485 1.185 ;
    END
  END q
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 11.995 1.015 12.325 1.185 ;
        RECT 15.235 1.015 15.565 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 3.435 0.085 3.605 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 12.075 0.085 12.245 1.015 ;
        RECT 15.315 0.085 15.485 1.015 ;
        RECT 0.000 -0.085 15.980 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
        RECT 10.965 -0.085 11.135 0.085 ;
        RECT 11.305 -0.085 11.475 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 11.985 -0.085 12.155 0.085 ;
        RECT 12.325 -0.085 12.495 0.085 ;
        RECT 12.665 -0.085 12.835 0.085 ;
        RECT 13.005 -0.085 13.175 0.085 ;
        RECT 13.345 -0.085 13.515 0.085 ;
        RECT 13.685 -0.085 13.855 0.085 ;
        RECT 14.025 -0.085 14.195 0.085 ;
        RECT 14.365 -0.085 14.535 0.085 ;
        RECT 14.705 -0.085 14.875 0.085 ;
        RECT 15.045 -0.085 15.215 0.085 ;
        RECT 15.385 -0.085 15.555 0.085 ;
        RECT 15.725 -0.085 15.895 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 15.980 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 15.980 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 12.075 3.055 12.245 3.995 ;
        RECT 15.315 3.055 15.485 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
        RECT 11.995 2.885 12.325 3.055 ;
        RECT 15.235 2.885 15.565 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
        RECT 10.965 3.995 11.135 4.165 ;
        RECT 11.305 3.995 11.475 4.165 ;
        RECT 11.645 3.995 11.815 4.165 ;
        RECT 11.985 3.995 12.155 4.165 ;
        RECT 12.325 3.995 12.495 4.165 ;
        RECT 12.665 3.995 12.835 4.165 ;
        RECT 13.005 3.995 13.175 4.165 ;
        RECT 13.345 3.995 13.515 4.165 ;
        RECT 13.685 3.995 13.855 4.165 ;
        RECT 14.025 3.995 14.195 4.165 ;
        RECT 14.365 3.995 14.535 4.165 ;
        RECT 14.705 3.995 14.875 4.165 ;
        RECT 15.045 3.995 15.215 4.165 ;
        RECT 15.385 3.995 15.555 4.165 ;
        RECT 15.725 3.995 15.895 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 15.980 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 16.160 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 15.675 1.395 ;
        RECT 0.005 0.485 2.715 0.715 ;
        RECT 7.565 0.710 9.195 0.715 ;
        RECT 11.885 0.485 15.675 0.715 ;
      LAYER li1 ;
        RECT 2.275 2.545 3.145 2.715 ;
        RECT 1.195 1.595 4.225 1.765 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 9.835 2.545 10.165 2.715 ;
        RECT 9.915 2.445 10.085 2.545 ;
        RECT 9.915 2.275 12.865 2.445 ;
        RECT 9.915 1.765 10.085 2.275 ;
        RECT 9.915 1.595 12.865 1.765 ;
        RECT 9.915 1.185 10.085 1.595 ;
        RECT 9.835 1.015 10.165 1.185 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 5.595 2.445 5.765 2.885 ;
        RECT 5.515 2.275 5.845 2.445 ;
        RECT 5.515 1.595 8.545 1.765 ;
        RECT 5.595 1.185 5.765 1.595 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 9.375 3.605 10.705 3.775 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 0.195 2.445 0.365 2.545 ;
        RECT 0.195 2.275 4.225 2.445 ;
        RECT 0.195 1.185 0.365 2.275 ;
        RECT 3.975 2.105 4.145 2.275 ;
        RECT 9.375 2.105 9.545 3.605 ;
        RECT 3.975 1.935 9.545 2.105 ;
        RECT 9.375 1.765 9.545 1.935 ;
        RECT 9.295 1.595 9.625 1.765 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 0.195 0.475 0.365 1.015 ;
        RECT 0.115 0.305 0.445 0.475 ;
        RECT 8.755 2.885 9.085 3.055 ;
        RECT 8.835 2.715 9.005 2.885 ;
        RECT 7.135 2.545 9.005 2.715 ;
        RECT 8.755 1.015 9.085 1.185 ;
        RECT 8.835 0.475 9.005 1.015 ;
        RECT 8.755 0.305 9.085 0.475 ;
        RECT 13.075 3.605 13.405 3.775 ;
        RECT 13.155 2.715 13.325 3.605 ;
        RECT 13.075 2.545 13.405 2.715 ;
        RECT 13.155 1.185 13.325 2.545 ;
        RECT 13.075 1.015 13.405 1.185 ;
        RECT 13.155 0.475 13.325 1.015 ;
        RECT 13.075 0.305 13.405 0.475 ;
  END
END DFQD1_3

#--------EOF---------

MACRO INVD1
  CLASS CORE ;
  FOREIGN INVD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.040 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 0.195 1.185 0.365 2.545 ;
        RECT 0.115 1.015 0.445 1.185 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 0.000 -0.085 2.040 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 2.040 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 2.040 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 2.040 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 2.220 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 1.635 1.395 ;
  END
END INVD1

#--------EOF---------

MACRO INVD1_1
  CLASS CORE ;
  FOREIGN INVD1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.040 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 0.195 1.185 0.365 2.545 ;
        RECT 0.115 1.015 0.445 1.185 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 0.000 -0.085 2.040 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 2.040 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 2.040 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 2.040 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 2.220 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 1.635 1.395 ;
  END
END INVD1_1

#--------EOF---------

MACRO INVD1_2
  CLASS CORE ;
  FOREIGN INVD1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.040 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 0.195 1.185 0.365 2.545 ;
        RECT 0.115 1.015 0.445 1.185 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 0.000 -0.085 2.040 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 2.040 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 2.040 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 2.040 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 2.220 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 1.635 1.395 ;
  END
END INVD1_2

#--------EOF---------

MACRO INVD1_3
  CLASS CORE ;
  FOREIGN INVD1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.040 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 0.195 1.185 0.365 2.545 ;
        RECT 0.115 1.015 0.445 1.185 ;
    END
  END z
  PIN i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END i
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 0.000 -0.085 2.040 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 2.040 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 2.040 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 2.040 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 2.220 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 1.635 1.395 ;
  END
END INVD1_3

#--------EOF---------

MACRO LNQD1
  CLASS CORE ;
  FOREIGN LNQD1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.880 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.105 0.905 2.445 ;
        RECT 0.655 1.935 0.985 2.105 ;
    END
  END en
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 9.835 2.545 10.165 2.715 ;
        RECT 9.915 1.185 10.085 2.545 ;
        RECT 9.835 1.015 10.165 1.185 ;
    END
  END q
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.177750 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END d
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 8.755 1.015 9.085 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 8.835 0.085 9.005 1.015 ;
        RECT 0.000 -0.085 10.880 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 10.880 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 10.880 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 8.835 3.055 9.005 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 8.755 2.885 9.085 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 10.880 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 11.060 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 10.275 1.395 ;
        RECT 1.085 0.700 3.795 0.715 ;
        RECT 8.645 0.485 10.275 0.715 ;
      LAYER li1 ;
        RECT 0.115 3.605 0.445 3.775 ;
        RECT 0.195 3.055 0.365 3.605 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 0.195 1.765 0.365 2.885 ;
        RECT 2.895 2.545 3.685 2.715 ;
        RECT 4.435 2.545 5.845 2.715 ;
        RECT 2.895 2.445 3.065 2.545 ;
        RECT 2.895 2.275 5.845 2.445 ;
        RECT 0.195 1.595 2.605 1.765 ;
        RECT 2.895 1.185 3.065 2.275 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.895 1.015 3.685 1.185 ;
        RECT 0.195 0.475 0.365 1.015 ;
        RECT 0.115 0.305 0.445 0.475 ;
        RECT 6.595 2.885 6.925 3.055 ;
        RECT 6.675 1.765 6.845 2.885 ;
        RECT 3.895 1.595 6.845 1.765 ;
        RECT 6.675 1.185 6.845 1.595 ;
        RECT 6.595 1.015 6.925 1.185 ;
        RECT 7.675 3.605 8.005 3.775 ;
        RECT 7.755 3.055 7.925 3.605 ;
        RECT 7.675 2.885 8.005 3.055 ;
        RECT 7.755 1.185 7.925 2.885 ;
        RECT 7.675 1.015 8.005 1.185 ;
  END
END LNQD1

#--------EOF---------

MACRO LNQD1_1
  CLASS CORE ;
  FOREIGN LNQD1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.880 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END en
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 9.835 2.545 10.165 2.715 ;
        RECT 9.915 1.185 10.085 2.545 ;
        RECT 9.835 1.015 10.165 1.185 ;
    END
  END q
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.177750 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END d
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 8.755 1.015 9.085 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 8.835 0.085 9.005 1.015 ;
        RECT 0.000 -0.085 10.880 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 10.880 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 10.880 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 8.835 3.055 9.005 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 8.755 2.885 9.085 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 10.880 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 11.060 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 10.275 1.395 ;
        RECT 1.085 0.700 3.795 0.715 ;
        RECT 8.645 0.485 10.275 0.715 ;
      LAYER li1 ;
        RECT 0.115 3.605 0.445 3.775 ;
        RECT 0.195 3.055 0.365 3.605 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 0.195 1.185 0.365 2.885 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 0.195 0.475 0.365 1.015 ;
        RECT 0.115 0.305 0.445 0.475 ;
        RECT 3.355 2.545 5.845 2.715 ;
        RECT 3.435 1.185 3.605 2.545 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 7.675 2.885 8.005 3.055 ;
        RECT 3.895 2.275 4.225 2.445 ;
        RECT 3.975 1.765 4.145 2.275 ;
        RECT 7.755 1.765 7.925 2.885 ;
        RECT 3.895 1.595 7.925 1.765 ;
        RECT 7.755 1.185 7.925 1.595 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 6.135 2.885 6.925 3.055 ;
        RECT 6.135 2.445 6.305 2.885 ;
        RECT 6.055 2.275 6.385 2.445 ;
        RECT 6.595 1.015 6.925 1.185 ;
        RECT 6.675 0.475 6.845 1.015 ;
        RECT 6.595 0.305 6.925 0.475 ;
  END
END LNQD1_1

#--------EOF---------

MACRO LNQD1_2
  CLASS CORE ;
  FOREIGN LNQD1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.900 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.105 0.905 2.445 ;
        RECT 0.655 1.935 0.985 2.105 ;
    END
  END en
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 9.295 2.545 10.165 2.715 ;
        RECT 9.295 1.015 10.165 1.185 ;
    END
  END q
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.177750 ;
    PORT
      LAYER li1 ;
        RECT 3.975 1.765 4.145 2.105 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END d
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 10.915 1.015 11.245 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 3.435 0.085 3.605 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 10.995 0.085 11.165 1.015 ;
        RECT 0.000 -0.085 11.900 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
        RECT 10.965 -0.085 11.135 0.085 ;
        RECT 11.305 -0.085 11.475 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 11.900 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 11.900 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 10.995 3.055 11.165 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
        RECT 10.915 2.885 11.245 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
        RECT 10.965 3.995 11.135 4.165 ;
        RECT 11.305 3.995 11.475 4.165 ;
        RECT 11.645 3.995 11.815 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 11.900 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 12.080 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 11.355 1.395 ;
        RECT 3.245 0.700 5.955 0.715 ;
        RECT 9.725 0.485 11.355 0.715 ;
      LAYER li1 ;
        RECT 0.115 3.605 0.445 3.775 ;
        RECT 0.195 3.055 0.365 3.605 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 0.195 2.715 0.365 2.885 ;
        RECT 0.195 2.545 2.065 2.715 ;
        RECT 0.195 1.765 0.365 2.545 ;
        RECT 0.195 1.595 2.065 1.765 ;
        RECT 0.195 1.185 0.365 1.595 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 5.515 2.545 8.545 2.715 ;
        RECT 5.595 1.765 5.765 2.545 ;
        RECT 5.595 1.595 10.705 1.765 ;
        RECT 5.595 1.185 5.765 1.595 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 2.355 2.445 2.525 2.885 ;
        RECT 2.355 2.275 5.305 2.445 ;
        RECT 2.355 1.185 2.525 2.275 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 5.055 0.475 5.225 2.275 ;
        RECT 5.055 0.305 6.385 0.475 ;
        RECT 8.755 2.885 9.085 3.055 ;
        RECT 8.835 2.715 9.005 2.885 ;
        RECT 8.755 2.545 9.085 2.715 ;
        RECT 8.755 1.015 9.085 1.185 ;
        RECT 8.835 0.475 9.005 1.015 ;
        RECT 8.755 0.305 9.085 0.475 ;
  END
END LNQD1_2

#--------EOF---------

MACRO LNQD1_3
  CLASS CORE ;
  FOREIGN LNQD1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.900 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.138000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END en
  PIN q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 9.295 2.545 10.165 2.715 ;
        RECT 9.295 1.015 10.165 1.185 ;
    END
  END q
  PIN d
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.177750 ;
    PORT
      LAYER li1 ;
        RECT 3.975 1.765 4.145 2.105 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END d
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 10.915 1.015 11.245 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 3.435 0.085 3.605 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 10.995 0.085 11.165 1.015 ;
        RECT 0.000 -0.085 11.900 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
        RECT 10.965 -0.085 11.135 0.085 ;
        RECT 11.305 -0.085 11.475 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 11.900 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 11.900 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 10.995 3.055 11.165 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
        RECT 10.915 2.885 11.245 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
        RECT 10.965 3.995 11.135 4.165 ;
        RECT 11.305 3.995 11.475 4.165 ;
        RECT 11.645 3.995 11.815 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 11.900 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 12.080 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 11.355 1.395 ;
        RECT 3.245 0.700 5.955 0.715 ;
        RECT 9.725 0.485 11.355 0.715 ;
      LAYER li1 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 2.355 2.715 2.525 2.885 ;
        RECT 0.655 2.545 2.525 2.715 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 2.355 0.475 2.525 1.015 ;
        RECT 2.275 0.305 2.605 0.475 ;
        RECT 5.515 2.545 8.545 2.715 ;
        RECT 6.135 1.765 6.305 2.545 ;
        RECT 6.135 1.595 10.705 1.765 ;
        RECT 6.135 1.185 6.305 1.595 ;
        RECT 5.515 1.015 6.305 1.185 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 0.195 2.445 0.365 2.885 ;
        RECT 0.195 2.275 5.305 2.445 ;
        RECT 0.195 1.185 0.365 2.275 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 8.755 2.885 9.085 3.055 ;
        RECT 8.835 2.715 9.005 2.885 ;
        RECT 8.755 2.545 9.085 2.715 ;
        RECT 8.755 1.015 9.085 1.185 ;
        RECT 8.835 0.475 9.005 1.015 ;
        RECT 8.755 0.305 9.085 0.475 ;
  END
END LNQD1_3

#--------EOF---------

MACRO MUX2D1
  CLASS CORE ;
  FOREIGN MUX2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 0.735 0.475 0.905 1.185 ;
        RECT 0.655 0.305 0.985 0.475 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.735 1.595 2.065 1.765 ;
        RECT 1.815 1.015 1.985 1.595 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.194250 ;
    PORT
      LAYER li1 ;
        RECT 2.815 1.595 3.145 1.765 ;
        RECT 2.895 1.015 3.065 1.595 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.823500 ;
    PORT
      LAYER li1 ;
        RECT 7.675 2.545 8.005 2.715 ;
        RECT 7.755 1.185 7.925 2.545 ;
        RECT 7.675 1.015 8.005 1.185 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 6.595 1.015 6.925 1.185 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 6.675 0.085 6.845 1.015 ;
        RECT 0.000 -0.085 8.500 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.500 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 8.500 4.165 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 6.675 3.055 6.845 3.995 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 6.595 2.885 6.925 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 8.500 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 8.680 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 8.115 1.395 ;
        RECT 1.085 0.665 3.795 0.715 ;
        RECT 1.085 0.485 2.715 0.665 ;
        RECT 6.485 0.485 8.115 0.715 ;
      LAYER li1 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 1.275 2.445 1.445 2.885 ;
        RECT 1.195 2.275 1.525 2.445 ;
        RECT 1.195 1.595 1.525 1.765 ;
        RECT 1.275 1.185 1.445 1.595 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 0.115 3.605 0.445 3.775 ;
        RECT 4.435 3.605 4.765 3.775 ;
        RECT 0.195 3.055 0.365 3.605 ;
        RECT 4.515 3.055 4.685 3.605 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
        RECT 0.195 1.185 0.365 2.885 ;
        RECT 4.515 1.595 5.845 1.765 ;
        RECT 4.515 1.185 4.685 1.595 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 3.355 2.545 4.145 2.715 ;
        RECT 3.975 1.185 4.145 2.545 ;
        RECT 3.355 1.015 4.145 1.185 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 5.595 2.715 5.765 2.885 ;
        RECT 4.515 2.545 6.305 2.715 ;
        RECT 4.515 2.105 4.685 2.545 ;
        RECT 0.655 1.935 3.685 2.105 ;
        RECT 4.435 1.935 4.765 2.105 ;
        RECT 6.135 1.185 6.305 2.545 ;
        RECT 5.515 1.015 6.305 1.185 ;
  END
END MUX2D1

#--------EOF---------

MACRO MUX2D1_1
  CLASS CORE ;
  FOREIGN MUX2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.105 3.065 2.445 ;
        RECT 2.815 1.935 3.145 2.105 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.203250 ;
    PORT
      LAYER li1 ;
        RECT 3.895 2.275 4.225 2.445 ;
        RECT 3.975 1.765 4.145 2.275 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.823500 ;
    PORT
      LAYER li1 ;
        RECT 6.595 2.545 6.925 2.715 ;
        RECT 6.675 1.185 6.845 2.545 ;
        RECT 6.595 1.015 6.925 1.185 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 0.000 -0.085 8.500 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.500 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 8.500 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 8.500 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 8.680 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 8.115 1.395 ;
        RECT 0.005 0.485 1.635 0.715 ;
        RECT 3.245 0.665 4.875 0.715 ;
        RECT 6.485 0.485 8.115 0.715 ;
      LAYER li1 ;
        RECT 1.195 2.545 1.525 2.715 ;
        RECT 1.275 1.185 1.445 2.545 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 2.275 3.605 2.605 3.775 ;
        RECT 2.355 3.055 2.525 3.605 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 2.355 1.185 2.525 2.885 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 3.435 1.185 3.605 2.885 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 1.735 2.545 2.065 2.715 ;
        RECT 1.815 0.475 1.985 2.545 ;
        RECT 5.595 1.185 5.765 2.885 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 5.595 0.475 5.765 1.015 ;
        RECT 1.815 0.305 3.145 0.475 ;
        RECT 5.515 0.305 5.845 0.475 ;
  END
END MUX2D1_1

#--------EOF---------

MACRO MUX2D1_2
  CLASS CORE ;
  FOREIGN MUX2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 1.735 1.935 4.145 2.105 ;
        RECT 3.975 1.765 4.145 1.935 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.815 1.595 3.145 1.765 ;
        RECT 2.895 1.015 3.065 1.595 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.194250 ;
    PORT
      LAYER li1 ;
        RECT 1.735 1.595 2.065 1.765 ;
        RECT 1.815 1.015 1.985 1.595 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.823500 ;
    PORT
      LAYER li1 ;
        RECT 7.675 2.545 8.005 2.715 ;
        RECT 7.755 1.185 7.925 2.545 ;
        RECT 7.675 1.015 8.005 1.185 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 6.595 1.015 6.925 1.185 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 6.675 0.085 6.845 1.015 ;
        RECT 0.000 -0.085 8.500 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.500 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 8.500 4.165 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 6.675 3.055 6.845 3.995 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 6.595 2.885 6.925 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 8.500 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 8.680 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 8.115 1.395 ;
        RECT 1.085 0.665 3.795 0.715 ;
        RECT 2.165 0.485 3.795 0.665 ;
        RECT 6.485 0.485 8.115 0.715 ;
      LAYER li1 ;
        RECT 3.355 2.545 3.685 2.715 ;
        RECT 3.435 2.445 3.605 2.545 ;
        RECT 3.355 2.275 3.685 2.445 ;
        RECT 3.355 1.595 3.685 1.765 ;
        RECT 3.435 1.185 3.605 1.595 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 0.115 3.605 0.445 3.775 ;
        RECT 4.435 3.605 4.765 3.775 ;
        RECT 0.195 3.055 0.365 3.605 ;
        RECT 4.515 3.055 4.685 3.605 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
        RECT 0.195 1.185 0.365 2.885 ;
        RECT 4.515 1.185 4.685 2.885 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 5.595 2.715 5.765 2.885 ;
        RECT 5.515 2.545 5.845 2.715 ;
        RECT 5.595 1.185 5.765 2.545 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 5.595 0.475 5.765 1.015 ;
        RECT 5.515 0.305 5.845 0.475 ;
  END
END MUX2D1_2

#--------EOF---------

MACRO MUX2D1_3
  CLASS CORE ;
  FOREIGN MUX2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN s
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 2.355 2.105 2.525 2.445 ;
        RECT 2.275 1.935 2.605 2.105 ;
    END
  END s
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.256500 ;
    PORT
      LAYER li1 ;
        RECT 3.895 2.275 4.225 2.445 ;
        RECT 3.975 1.765 4.145 2.275 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END i1
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.194250 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END i0
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.823500 ;
    PORT
      LAYER li1 ;
        RECT 6.595 2.545 6.925 2.715 ;
        RECT 6.675 1.185 6.845 2.545 ;
        RECT 6.595 1.015 6.925 1.185 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 0.000 -0.085 8.500 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.500 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 8.500 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 8.500 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 8.680 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 8.115 1.395 ;
        RECT 0.005 0.665 1.635 0.715 ;
        RECT 3.245 0.485 4.875 0.715 ;
        RECT 6.485 0.485 8.115 0.715 ;
      LAYER li1 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 3.435 1.185 3.605 2.885 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 2.815 3.605 3.145 3.775 ;
        RECT 2.895 3.055 3.065 3.605 ;
        RECT 2.275 2.885 3.065 3.055 ;
        RECT 2.895 1.185 3.065 2.885 ;
        RECT 2.275 1.015 3.065 1.185 ;
        RECT 1.195 2.545 1.525 2.715 ;
        RECT 1.275 1.185 1.445 2.545 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 1.815 2.545 2.605 2.715 ;
        RECT 1.815 1.765 1.985 2.545 ;
        RECT 1.735 1.595 2.065 1.765 ;
        RECT 5.595 1.185 5.765 2.885 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 5.595 0.475 5.765 1.015 ;
        RECT 5.515 0.305 5.845 0.475 ;
  END
END MUX2D1_3

#--------EOF---------

MACRO ND2D1
  CLASS CORE ;
  FOREIGN ND2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.060 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.326500 ;
    PORT
      LAYER li1 ;
        RECT 1.195 2.545 1.525 2.715 ;
        RECT 1.275 1.765 1.445 2.545 ;
        RECT 1.275 1.595 2.525 1.765 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 2.275 1.015 2.605 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 0.000 -0.085 3.060 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.060 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 3.060 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 2.275 2.885 2.605 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 3.060 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 3.240 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 2.715 1.395 ;
  END
END ND2D1

#--------EOF---------

MACRO ND2D1_1
  CLASS CORE ;
  FOREIGN ND2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.060 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.326500 ;
    PORT
      LAYER li1 ;
        RECT 1.195 2.545 1.525 2.715 ;
        RECT 1.275 2.445 1.445 2.545 ;
        RECT 0.195 2.275 1.445 2.445 ;
        RECT 0.195 1.185 0.365 2.275 ;
        RECT 0.115 1.015 0.445 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 0.000 -0.085 3.060 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.060 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 3.060 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 2.275 2.885 2.605 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 3.060 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 3.240 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 2.715 1.395 ;
  END
END ND2D1_1

#--------EOF---------

MACRO ND2D1_2
  CLASS CORE ;
  FOREIGN ND2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.060 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.616500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.545 2.605 2.715 ;
        RECT 1.815 1.185 1.985 2.545 ;
        RECT 1.815 1.015 2.605 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.275 1.765 1.445 2.105 ;
        RECT 1.195 1.595 1.525 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 0.000 -0.085 3.060 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.060 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 3.060 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 3.060 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 3.240 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 2.715 1.395 ;
  END
END ND2D1_2

#--------EOF---------

MACRO ND2D1_3
  CLASS CORE ;
  FOREIGN ND2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.060 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.616500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.545 2.605 2.715 ;
        RECT 0.195 1.185 0.365 2.545 ;
        RECT 0.115 1.015 0.445 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 0.000 -0.085 3.060 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.060 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 3.060 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 3.060 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 3.240 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 2.715 1.395 ;
  END
END ND2D1_3

#--------EOF---------

MACRO ND3D1
  CLASS CORE ;
  FOREIGN ND3D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.936500 ;
    PORT
      LAYER li1 ;
        RECT 1.195 2.545 3.685 2.715 ;
        RECT 1.275 1.765 1.445 2.545 ;
        RECT 1.275 1.595 2.525 1.765 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 2.275 1.015 2.605 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.975 1.765 4.145 2.105 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 0.000 -0.085 5.440 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 5.440 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 5.440 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 5.620 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 4.875 1.395 ;
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 0.195 0.475 0.365 1.015 ;
        RECT 3.435 0.475 3.605 1.015 ;
        RECT 0.195 0.305 3.605 0.475 ;
  END
END ND3D1

#--------EOF---------

MACRO ND3D1_1
  CLASS CORE ;
  FOREIGN ND3D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.080 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.936500 ;
    PORT
      LAYER li1 ;
        RECT 1.195 2.545 3.685 2.715 ;
        RECT 3.435 1.185 3.605 2.545 ;
        RECT 3.355 1.015 3.685 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 1.765 3.065 2.105 ;
        RECT 2.815 1.595 3.145 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 0.000 -0.085 4.080 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.080 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 4.080 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 2.275 2.885 2.605 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 4.080 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 4.260 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 3.795 1.395 ;
  END
END ND3D1_1

#--------EOF---------

MACRO ND3D1_2
  CLASS CORE ;
  FOREIGN ND3D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.936500 ;
    PORT
      LAYER li1 ;
        RECT 1.195 2.545 3.685 2.715 ;
        RECT 1.815 2.105 1.985 2.545 ;
        RECT 1.815 1.935 3.065 2.105 ;
        RECT 2.895 1.185 3.065 1.935 ;
        RECT 2.895 1.015 3.685 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.975 2.105 4.145 2.445 ;
        RECT 3.895 1.935 4.225 2.105 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.275 1.765 1.445 2.105 ;
        RECT 1.195 1.595 1.525 1.765 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 0.000 -0.085 5.440 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 5.440 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 5.440 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 5.620 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 4.875 1.395 ;
      LAYER li1 ;
        RECT 1.815 1.595 2.605 1.765 ;
        RECT 3.355 1.595 4.685 1.765 ;
        RECT 1.815 1.185 1.985 1.595 ;
        RECT 4.515 1.185 4.685 1.595 ;
        RECT 0.115 1.015 1.985 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
  END
END ND3D1_2

#--------EOF---------

MACRO ND3D1_3
  CLASS CORE ;
  FOREIGN ND3D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.080 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.936500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.545 2.605 2.715 ;
        RECT 0.195 1.185 0.365 2.545 ;
        RECT 0.115 1.015 0.445 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 1.765 3.065 2.105 ;
        RECT 2.815 1.595 3.145 1.765 ;
    END
  END a3
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 3.435 0.085 3.605 1.015 ;
        RECT 0.000 -0.085 4.080 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.080 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 4.080 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 3.355 2.885 3.685 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 4.080 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 4.260 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 3.795 1.395 ;
  END
END ND3D1_3

#--------EOF---------

MACRO ND4D1
  CLASS CORE ;
  FOREIGN ND4D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 5.055 1.765 5.225 2.105 ;
        RECT 4.975 1.595 5.305 1.765 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.975 1.765 4.145 2.105 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END a3
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.256500 ;
    PORT
      LAYER li1 ;
        RECT 1.195 2.545 4.765 2.715 ;
        RECT 1.275 1.185 1.445 2.545 ;
        RECT 1.275 1.015 2.605 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 0.000 -0.085 6.460 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.460 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 6.460 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 6.460 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 6.640 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 5.955 1.395 ;
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 0.195 0.475 0.365 1.015 ;
        RECT 3.435 0.475 3.605 1.015 ;
        RECT 0.195 0.305 3.605 0.475 ;
  END
END ND4D1

#--------EOF---------

MACRO ND4D1_1
  CLASS CORE ;
  FOREIGN ND4D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a2
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 5.055 1.765 5.225 2.105 ;
        RECT 4.975 1.595 5.305 1.765 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a3
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.546500 ;
    PORT
      LAYER li1 ;
        RECT 1.195 2.545 4.765 2.715 ;
        RECT 2.895 1.185 3.065 2.545 ;
        RECT 2.895 1.015 3.685 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.355 1.765 2.525 2.105 ;
        RECT 2.275 1.595 2.605 1.765 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 0.000 -0.085 6.460 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.460 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 6.460 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 6.460 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 6.640 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 5.955 1.395 ;
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 0.195 0.475 0.365 1.015 ;
        RECT 4.515 0.475 4.685 1.015 ;
        RECT 0.195 0.305 4.685 0.475 ;
  END
END ND4D1_1

#--------EOF---------

MACRO ND4D1_2
  CLASS CORE ;
  FOREIGN ND4D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a3
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.546500 ;
    PORT
      LAYER li1 ;
        RECT 1.195 2.545 4.765 2.715 ;
        RECT 3.435 1.765 3.605 2.545 ;
        RECT 3.435 1.595 4.685 1.765 ;
        RECT 4.515 1.185 4.685 1.595 ;
        RECT 4.435 1.015 4.765 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 5.055 1.765 5.225 2.105 ;
        RECT 4.975 1.595 5.305 1.765 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 3.435 0.085 3.605 1.015 ;
        RECT 0.000 -0.085 6.460 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.460 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 6.460 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 6.460 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 6.640 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 5.955 1.395 ;
      LAYER li1 ;
        RECT 2.895 1.765 3.065 2.105 ;
        RECT 2.815 1.595 3.145 1.765 ;
        RECT 0.115 1.015 3.065 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 2.895 0.475 3.065 1.015 ;
        RECT 5.595 0.475 5.765 1.015 ;
        RECT 2.815 0.305 3.145 0.475 ;
        RECT 5.515 0.305 5.845 0.475 ;
  END
END ND4D1_2

#--------EOF---------

MACRO ND4D1_3
  CLASS CORE ;
  FOREIGN ND4D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.105 3.065 2.445 ;
        RECT 2.815 1.935 3.145 2.105 ;
    END
  END a2
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END a3
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.256500 ;
    PORT
      LAYER li1 ;
        RECT 1.195 2.545 1.525 2.715 ;
        RECT 3.355 2.545 3.685 2.715 ;
        RECT 1.275 1.765 1.445 2.545 ;
        RECT 3.435 1.765 3.605 2.545 ;
        RECT 1.275 1.595 4.685 1.765 ;
        RECT 4.515 1.185 4.685 1.595 ;
        RECT 4.435 1.015 4.765 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.975 2.105 4.145 2.445 ;
        RECT 3.895 1.935 4.225 2.105 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 0.000 -0.085 5.440 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 5.440 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 5.440 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 5.620 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 4.875 1.395 ;
  END
END ND4D1_3

#--------EOF---------

MACRO NR2D1
  CLASS CORE ;
  FOREIGN NR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.060 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.214500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 0.195 1.765 0.365 2.545 ;
        RECT 0.195 1.595 1.445 1.765 ;
        RECT 1.275 1.185 1.445 1.595 ;
        RECT 1.195 1.015 1.525 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.105 0.905 2.445 ;
        RECT 0.655 1.935 0.985 2.105 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 0.000 -0.085 3.060 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.060 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 3.060 4.165 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 2.275 2.885 2.605 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 3.060 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 3.240 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 2.715 1.395 ;
  END
END NR2D1

#--------EOF---------

MACRO NR2D1_1
  CLASS CORE ;
  FOREIGN NR2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.060 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.214500 ;
    PORT
      LAYER li1 ;
        RECT 2.275 2.545 2.605 2.715 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 1.275 2.275 2.525 2.445 ;
        RECT 1.275 1.185 1.445 2.275 ;
        RECT 1.195 1.015 1.525 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 0.000 -0.085 3.060 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.060 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 3.060 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 3.060 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 3.240 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 2.715 1.395 ;
  END
END NR2D1_1

#--------EOF---------

MACRO NR2D1_2
  CLASS CORE ;
  FOREIGN NR2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.060 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.403000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 0.195 1.765 0.365 2.545 ;
        RECT 0.195 1.595 2.525 1.765 ;
        RECT 0.195 1.185 0.365 1.595 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.105 0.905 2.445 ;
        RECT 0.655 1.935 0.985 2.105 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 0.000 -0.085 3.060 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.060 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 3.060 4.165 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 2.275 2.885 2.605 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 3.060 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 3.240 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 2.715 1.395 ;
  END
END NR2D1_2

#--------EOF---------

MACRO NR2D1_3
  CLASS CORE ;
  FOREIGN NR2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.060 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.403000 ;
    PORT
      LAYER li1 ;
        RECT 0.195 2.545 2.605 2.715 ;
        RECT 0.195 1.185 0.365 2.545 ;
        RECT 2.355 1.185 2.525 2.545 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 0.000 -0.085 3.060 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 3.060 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 3.060 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 3.060 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 3.240 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 2.715 1.395 ;
  END
END NR2D1_3

#--------EOF---------

MACRO NR3D1
  CLASS CORE ;
  FOREIGN NR3D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.880 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.146500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.885 5.225 3.055 ;
        RECT 5.055 2.715 5.225 2.885 ;
        RECT 1.195 2.545 1.525 2.715 ;
        RECT 5.055 2.545 9.085 2.715 ;
        RECT 1.275 1.765 1.445 2.545 ;
        RECT 1.275 1.595 3.605 1.765 ;
        RECT 1.275 1.185 1.445 1.595 ;
        RECT 3.435 1.185 3.605 1.595 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.397500 ;
    ANTENNADIFFAREA 1.215500 ;
    PORT
      LAYER li1 ;
        RECT 7.135 3.605 7.465 3.775 ;
        RECT 9.835 3.605 10.165 3.775 ;
        RECT 7.215 3.055 7.385 3.605 ;
        RECT 9.915 3.055 10.085 3.605 ;
        RECT 6.595 2.885 7.385 3.055 ;
        RECT 9.835 2.885 10.165 3.055 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 0.195 1.765 0.365 2.105 ;
        RECT 1.735 1.935 2.065 2.105 ;
        RECT 0.115 1.595 0.445 1.765 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.415500 ;
    PORT
      LAYER li1 ;
        RECT 2.815 2.275 9.625 2.445 ;
        RECT 3.975 1.765 4.145 2.275 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.397500 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.935 0.985 2.105 ;
        RECT 0.735 0.475 0.905 1.935 ;
        RECT 0.735 0.305 2.065 0.475 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 6.595 1.015 6.925 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 8.755 1.015 9.085 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 6.675 0.085 6.845 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 8.835 0.085 9.005 1.015 ;
        RECT 0.000 -0.085 10.880 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 10.880 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 10.880 4.165 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 10.880 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 11.060 4.405 ;
      LAYER pwell ;
        RECT 0.005 1.375 3.795 1.395 ;
        RECT 0.005 0.825 9.195 1.375 ;
        RECT 0.005 0.485 3.795 0.825 ;
      LAYER li1 ;
        RECT 3.355 2.545 4.765 2.715 ;
  END
END NR3D1

#--------EOF---------

MACRO NR3D1_1
  CLASS CORE ;
  FOREIGN NR3D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.900 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.146500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.885 3.685 3.055 ;
        RECT 1.195 2.545 1.525 2.715 ;
        RECT 1.275 1.765 1.445 2.545 ;
        RECT 1.275 1.595 3.605 1.765 ;
        RECT 1.275 1.185 1.445 1.595 ;
        RECT 3.435 1.185 3.605 1.595 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.397500 ;
    ANTENNADIFFAREA 1.215500 ;
    PORT
      LAYER li1 ;
        RECT 8.215 3.605 8.545 3.775 ;
        RECT 10.915 3.605 11.245 3.775 ;
        RECT 8.295 3.055 8.465 3.605 ;
        RECT 10.995 3.055 11.165 3.605 ;
        RECT 7.675 2.885 8.465 3.055 ;
        RECT 10.915 2.885 11.245 3.055 ;
        RECT 3.435 2.105 3.605 2.445 ;
        RECT 3.355 1.935 3.685 2.105 ;
        RECT 1.735 0.305 2.065 0.475 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.415500 ;
    PORT
      LAYER li1 ;
        RECT 3.895 2.275 10.705 2.445 ;
        RECT 3.975 1.765 4.145 2.275 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.397500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 6.595 1.015 6.925 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 8.755 1.015 9.085 1.185 ;
        RECT 9.835 1.015 10.165 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 6.675 0.085 6.845 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 8.835 0.085 9.005 1.015 ;
        RECT 9.915 0.085 10.085 1.015 ;
        RECT 0.000 -0.085 11.900 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
        RECT 10.965 -0.085 11.135 0.085 ;
        RECT 11.305 -0.085 11.475 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 11.900 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 11.900 4.165 ;
        RECT 6.675 3.055 6.845 3.995 ;
        RECT 8.835 3.055 9.005 3.995 ;
        RECT 6.595 2.885 6.925 3.055 ;
        RECT 8.755 2.885 9.085 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
        RECT 10.965 3.995 11.135 4.165 ;
        RECT 11.305 3.995 11.475 4.165 ;
        RECT 11.645 3.995 11.815 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 11.900 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 12.080 4.405 ;
      LAYER pwell ;
        RECT 0.005 1.375 4.875 1.395 ;
        RECT 0.005 0.825 10.275 1.375 ;
        RECT 0.005 0.485 4.875 0.825 ;
      LAYER li1 ;
        RECT 2.275 2.545 10.165 2.715 ;
        RECT 4.435 2.885 5.845 3.055 ;
  END
END NR3D1_1

#--------EOF---------

MACRO NR3D1_2
  CLASS CORE ;
  FOREIGN NR3D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.880 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.397500 ;
    ANTENNADIFFAREA 4.362000 ;
    PORT
      LAYER li1 ;
        RECT 3.435 3.605 4.685 3.775 ;
        RECT 4.975 3.605 5.305 3.775 ;
        RECT 8.755 3.605 9.085 3.775 ;
        RECT 3.435 3.055 3.605 3.605 ;
        RECT 4.515 3.055 4.685 3.605 ;
        RECT 5.055 3.055 5.225 3.605 ;
        RECT 8.835 3.055 9.005 3.605 ;
        RECT 0.115 2.885 5.225 3.055 ;
        RECT 8.755 2.885 9.085 3.055 ;
        RECT 1.195 2.545 1.525 2.715 ;
        RECT 1.275 2.445 1.445 2.545 ;
        RECT 0.195 2.275 1.985 2.445 ;
        RECT 0.195 1.765 0.365 2.275 ;
        RECT 1.195 1.935 1.525 2.105 ;
        RECT 0.195 1.595 2.525 1.765 ;
        RECT 0.195 1.185 0.365 1.595 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 0.655 0.305 0.985 0.475 ;
    END
  END zn
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.415500 ;
    PORT
      LAYER li1 ;
        RECT 2.815 2.275 9.625 2.445 ;
        RECT 2.895 1.765 3.065 2.275 ;
        RECT 2.815 1.595 3.145 1.765 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.414000 ;
    PORT
      LAYER li1 ;
        RECT 2.355 2.545 8.545 2.715 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 2.275 2.275 2.605 2.445 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 6.595 1.015 6.925 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 8.755 1.015 9.085 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 3.435 0.085 3.605 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 6.675 0.085 6.845 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 8.835 0.085 9.005 1.015 ;
        RECT 0.000 -0.085 10.880 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 10.880 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 10.880 4.165 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 10.880 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 11.060 4.405 ;
      LAYER pwell ;
        RECT 0.005 1.375 3.795 1.395 ;
        RECT 0.005 0.825 9.195 1.375 ;
        RECT 0.005 0.485 3.795 0.825 ;
  END
END NR3D1_2

#--------EOF---------

MACRO NR3D1_3
  CLASS CORE ;
  FOREIGN NR3D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.880 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.931000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 2.275 2.545 2.605 2.715 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 1.275 2.275 2.525 2.445 ;
        RECT 1.275 1.765 1.445 2.275 ;
        RECT 1.275 1.595 3.605 1.765 ;
        RECT 1.275 1.185 1.445 1.595 ;
        RECT 3.435 1.185 3.605 1.595 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
    END
  END zn
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.397500 ;
    ANTENNADIFFAREA 1.215500 ;
    PORT
      LAYER li1 ;
        RECT 7.135 3.605 7.465 3.775 ;
        RECT 9.835 3.605 10.165 3.775 ;
        RECT 7.215 3.055 7.385 3.605 ;
        RECT 9.915 3.055 10.085 3.605 ;
        RECT 6.595 2.885 7.385 3.055 ;
        RECT 9.835 2.885 10.165 3.055 ;
        RECT 3.975 1.765 4.145 2.105 ;
        RECT 3.895 1.595 4.225 1.765 ;
        RECT 2.815 0.305 3.145 0.475 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.819500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 3.605 2.065 3.775 ;
        RECT 0.735 0.475 0.905 3.605 ;
        RECT 3.355 2.275 9.625 2.445 ;
        RECT 0.655 0.305 0.985 0.475 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 6.595 1.015 6.925 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 8.755 1.015 9.085 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 6.675 0.085 6.845 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 8.835 0.085 9.005 1.015 ;
        RECT 0.000 -0.085 10.880 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 10.880 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 10.880 4.165 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 10.880 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 11.060 4.405 ;
      LAYER pwell ;
        RECT 0.005 1.375 3.795 1.395 ;
        RECT 0.005 0.825 9.195 1.375 ;
        RECT 0.005 0.485 3.795 0.825 ;
      LAYER li1 ;
        RECT 3.355 2.545 9.085 2.715 ;
  END
END NR3D1_3

#--------EOF---------

MACRO NR4D1
  CLASS CORE ;
  FOREIGN NR4D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.960 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.940500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.885 3.685 3.055 ;
        RECT 1.195 2.545 1.525 2.715 ;
        RECT 1.275 1.765 1.445 2.545 ;
        RECT 1.275 1.595 4.685 1.765 ;
        RECT 1.275 1.185 1.445 1.595 ;
        RECT 4.515 1.185 4.685 1.595 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
    END
  END zn
  PIN a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363750 ;
    ANTENNADIFFAREA 1.215500 ;
    PORT
      LAYER li1 ;
        RECT 9.295 3.605 9.625 3.775 ;
        RECT 14.155 3.605 14.485 3.775 ;
        RECT 9.375 3.055 9.545 3.605 ;
        RECT 14.235 3.055 14.405 3.605 ;
        RECT 8.755 2.885 9.545 3.055 ;
        RECT 14.155 2.885 14.485 3.055 ;
        RECT 5.055 1.765 5.225 2.105 ;
        RECT 4.975 1.595 5.305 1.765 ;
    END
  END a4
  PIN a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.388250 ;
    PORT
      LAYER li1 ;
        RECT 6.595 2.275 13.945 2.445 ;
    END
  END a3
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.380250 ;
    PORT
      LAYER li1 ;
        RECT 4.435 2.275 6.305 2.445 ;
        RECT 6.135 2.105 6.305 2.275 ;
        RECT 6.135 1.935 7.465 2.105 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.363750 ;
    PORT
      LAYER li1 ;
        RECT 0.655 1.935 0.985 2.105 ;
        RECT 0.735 0.475 0.905 1.935 ;
        RECT 0.735 0.305 2.065 0.475 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 6.595 1.015 6.925 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 8.755 1.015 9.085 1.185 ;
        RECT 9.835 1.015 10.165 1.185 ;
        RECT 10.915 1.015 11.245 1.185 ;
        RECT 11.995 1.015 12.325 1.185 ;
        RECT 13.075 1.015 13.405 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 3.435 0.085 3.605 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 6.675 0.085 6.845 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 8.835 0.085 9.005 1.015 ;
        RECT 9.915 0.085 10.085 1.015 ;
        RECT 10.995 0.085 11.165 1.015 ;
        RECT 12.075 0.085 12.245 1.015 ;
        RECT 13.155 0.085 13.325 1.015 ;
        RECT 0.000 -0.085 14.960 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
        RECT 8.585 -0.085 8.755 0.085 ;
        RECT 8.925 -0.085 9.095 0.085 ;
        RECT 9.265 -0.085 9.435 0.085 ;
        RECT 9.605 -0.085 9.775 0.085 ;
        RECT 9.945 -0.085 10.115 0.085 ;
        RECT 10.285 -0.085 10.455 0.085 ;
        RECT 10.625 -0.085 10.795 0.085 ;
        RECT 10.965 -0.085 11.135 0.085 ;
        RECT 11.305 -0.085 11.475 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 11.985 -0.085 12.155 0.085 ;
        RECT 12.325 -0.085 12.495 0.085 ;
        RECT 12.665 -0.085 12.835 0.085 ;
        RECT 13.005 -0.085 13.175 0.085 ;
        RECT 13.345 -0.085 13.515 0.085 ;
        RECT 13.685 -0.085 13.855 0.085 ;
        RECT 14.025 -0.085 14.195 0.085 ;
        RECT 14.365 -0.085 14.535 0.085 ;
        RECT 14.705 -0.085 14.875 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 14.960 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 14.960 4.165 ;
        RECT 9.915 3.055 10.085 3.995 ;
        RECT 12.075 3.055 12.245 3.995 ;
        RECT 9.835 2.885 10.165 3.055 ;
        RECT 11.995 2.885 12.325 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
        RECT 8.585 3.995 8.755 4.165 ;
        RECT 8.925 3.995 9.095 4.165 ;
        RECT 9.265 3.995 9.435 4.165 ;
        RECT 9.605 3.995 9.775 4.165 ;
        RECT 9.945 3.995 10.115 4.165 ;
        RECT 10.285 3.995 10.455 4.165 ;
        RECT 10.625 3.995 10.795 4.165 ;
        RECT 10.965 3.995 11.135 4.165 ;
        RECT 11.305 3.995 11.475 4.165 ;
        RECT 11.645 3.995 11.815 4.165 ;
        RECT 11.985 3.995 12.155 4.165 ;
        RECT 12.325 3.995 12.495 4.165 ;
        RECT 12.665 3.995 12.835 4.165 ;
        RECT 13.005 3.995 13.175 4.165 ;
        RECT 13.345 3.995 13.515 4.165 ;
        RECT 13.685 3.995 13.855 4.165 ;
        RECT 14.025 3.995 14.195 4.165 ;
        RECT 14.365 3.995 14.535 4.165 ;
        RECT 14.705 3.995 14.875 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 14.960 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 15.140 4.405 ;
      LAYER pwell ;
        RECT 0.005 1.375 5.955 1.395 ;
        RECT 0.005 0.825 13.515 1.375 ;
        RECT 0.005 0.710 5.955 0.825 ;
      LAYER li1 ;
        RECT 2.275 2.545 6.925 2.715 ;
        RECT 7.675 2.545 13.405 2.715 ;
  END
END NR4D1

#--------EOF---------

MACRO OA21D1
  CLASS CORE ;
  FOREIGN OA21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.105 3.065 2.445 ;
        RECT 2.815 1.935 3.145 2.105 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 4.435 2.545 4.765 2.715 ;
        RECT 4.515 1.185 4.685 2.545 ;
        RECT 4.435 1.015 4.765 1.185 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 0.000 -0.085 6.460 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.460 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 6.460 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 6.460 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 6.640 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 5.955 1.395 ;
      LAYER li1 ;
        RECT 1.195 2.545 3.605 2.715 ;
        RECT 3.435 1.765 3.605 2.545 ;
        RECT 3.355 1.595 4.145 1.765 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 2.355 0.475 2.525 1.015 ;
        RECT 3.975 0.475 4.145 1.595 ;
        RECT 2.355 0.305 4.145 0.475 ;
        RECT 1.275 1.595 3.065 1.765 ;
        RECT 1.275 1.185 1.445 1.595 ;
        RECT 2.895 1.185 3.065 1.595 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 2.895 1.015 3.685 1.185 ;
  END
END OA21D1

#--------EOF---------

MACRO OA21D1_1
  CLASS CORE ;
  FOREIGN OA21D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.105 0.905 2.445 ;
        RECT 0.655 1.935 0.985 2.105 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.105 3.065 2.445 ;
        RECT 2.815 1.935 3.145 2.105 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 4.435 2.545 4.765 2.715 ;
        RECT 4.515 1.185 4.685 2.545 ;
        RECT 4.435 1.015 4.765 1.185 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 3.435 0.085 3.605 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 0.000 -0.085 6.460 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.460 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 6.460 4.165 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 6.460 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 6.640 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 5.955 1.395 ;
      LAYER li1 ;
        RECT 3.435 3.605 5.305 3.775 ;
        RECT 3.435 3.055 3.605 3.605 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 1.275 2.545 3.685 2.715 ;
        RECT 0.195 1.765 0.365 2.545 ;
        RECT 1.275 1.765 1.445 2.545 ;
        RECT 0.195 1.595 4.225 1.765 ;
        RECT 1.275 1.185 1.445 1.595 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 0.195 0.475 0.365 1.015 ;
        RECT 2.355 0.475 2.525 1.015 ;
        RECT 0.195 0.305 2.525 0.475 ;
  END
END OA21D1_1

#--------EOF---------

MACRO OA21D1_2
  CLASS CORE ;
  FOREIGN OA21D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.975 1.765 4.145 2.105 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.002000 ;
    PORT
      LAYER li1 ;
        RECT 5.515 2.545 5.845 2.715 ;
        RECT 5.595 1.185 5.765 2.545 ;
        RECT 5.515 1.015 5.845 1.185 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 0.000 -0.085 6.460 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.460 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 6.460 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 6.460 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 6.640 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 5.955 1.395 ;
      LAYER li1 ;
        RECT 2.275 2.545 2.605 2.715 ;
        RECT 3.355 2.545 3.685 2.715 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 3.435 2.445 3.605 2.545 ;
        RECT 0.195 2.275 5.305 2.445 ;
        RECT 0.195 1.185 0.365 2.275 ;
        RECT 2.355 1.185 2.525 2.275 ;
        RECT 5.055 1.765 5.225 2.275 ;
        RECT 4.975 1.595 5.305 1.765 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 1.275 0.475 1.445 1.015 ;
        RECT 3.435 0.475 3.605 1.015 ;
        RECT 1.275 0.305 3.605 0.475 ;
  END
END OA21D1_2

#--------EOF---------

MACRO OA21D1_3
  CLASS CORE ;
  FOREIGN OA21D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.460 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END a2
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 2.105 3.065 2.445 ;
        RECT 2.815 1.935 3.145 2.105 ;
    END
  END a1
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END b
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 4.435 2.545 4.765 2.715 ;
        RECT 4.515 1.185 4.685 2.545 ;
        RECT 4.435 1.015 4.765 1.185 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 5.595 0.085 5.765 1.015 ;
        RECT 0.000 -0.085 6.460 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 6.460 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 6.460 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 5.595 3.055 5.765 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 5.515 2.885 5.845 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 6.460 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 6.640 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 5.955 1.395 ;
      LAYER li1 ;
        RECT 3.435 3.605 5.305 3.775 ;
        RECT 3.435 3.055 3.605 3.605 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 0.115 2.545 3.685 2.715 ;
        RECT 3.435 1.765 3.605 2.545 ;
        RECT 3.355 1.595 4.145 1.765 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 2.355 0.475 2.525 1.015 ;
        RECT 3.975 0.475 4.145 1.595 ;
        RECT 2.355 0.305 4.145 0.475 ;
        RECT 1.275 1.595 3.065 1.765 ;
        RECT 1.275 1.185 1.445 1.595 ;
        RECT 2.895 1.185 3.065 1.595 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 2.895 1.015 3.685 1.185 ;
  END
END OA21D1_3

#--------EOF---------

MACRO OAI21D1
  CLASS CORE ;
  FOREIGN OAI21D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.080 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.534500 ;
    PORT
      LAYER li1 ;
        RECT 1.195 2.545 1.525 2.715 ;
        RECT 1.275 1.765 1.445 2.545 ;
        RECT 1.275 1.595 2.525 1.765 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 2.275 1.015 2.605 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 1.765 3.065 2.105 ;
        RECT 2.815 1.595 3.145 1.765 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 0.000 -0.085 4.080 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.080 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 4.080 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 3.355 2.885 3.685 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 4.080 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 4.260 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 3.795 1.395 ;
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 1.275 0.475 1.445 1.015 ;
        RECT 3.435 0.475 3.605 1.015 ;
        RECT 1.275 0.305 3.605 0.475 ;
  END
END OAI21D1

#--------EOF---------

MACRO OAI21D1_1
  CLASS CORE ;
  FOREIGN OAI21D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.080 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.530000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 2.545 2.605 2.715 ;
        RECT 2.355 2.105 2.525 2.545 ;
        RECT 1.195 1.935 1.525 2.105 ;
        RECT 2.275 1.935 2.605 2.105 ;
        RECT 1.275 1.185 1.445 1.935 ;
        RECT 1.195 1.015 1.525 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.256500 ;
    PORT
      LAYER li1 ;
        RECT 1.735 2.275 2.065 2.445 ;
        RECT 1.815 1.765 1.985 2.275 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 1.765 3.065 2.105 ;
        RECT 2.815 1.595 3.145 1.765 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 3.435 0.085 3.605 1.015 ;
        RECT 0.000 -0.085 4.080 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.080 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 4.080 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 3.435 3.055 3.605 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 3.355 2.885 3.685 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 4.080 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 4.260 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 3.795 1.395 ;
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 0.195 0.475 0.365 1.015 ;
        RECT 2.355 0.475 2.525 1.015 ;
        RECT 0.195 0.305 2.525 0.475 ;
  END
END OAI21D1_1

#--------EOF---------

MACRO OAI21D1_2
  CLASS CORE ;
  FOREIGN OAI21D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.013000 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 2.895 2.545 3.685 2.715 ;
        RECT 0.195 1.185 0.365 2.545 ;
        RECT 2.895 1.185 3.065 2.545 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 3.065 1.185 ;
        RECT 0.195 0.475 0.365 1.015 ;
        RECT 2.355 0.475 2.525 1.015 ;
        RECT 0.195 0.305 2.525 0.475 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.975 1.765 4.145 2.105 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 0.000 -0.085 5.440 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 5.440 4.165 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 5.440 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 5.620 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 4.875 1.395 ;
      LAYER li1 ;
        RECT 1.275 1.595 2.605 1.765 ;
        RECT 3.355 1.595 3.685 1.765 ;
        RECT 1.275 1.185 1.445 1.595 ;
        RECT 3.435 1.185 3.605 1.595 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
  END
END OAI21D1_2

#--------EOF---------

MACRO OAI21D1_3
  CLASS CORE ;
  FOREIGN OAI21D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.013000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 2.545 3.685 2.715 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 0.195 2.275 2.525 2.445 ;
        RECT 0.195 1.185 0.365 2.275 ;
        RECT 2.355 1.185 2.525 2.275 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.975 1.765 4.145 2.105 ;
        RECT 3.895 1.595 4.225 1.765 ;
    END
  END b
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 0.000 -0.085 5.440 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 5.440 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 5.440 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 5.620 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 4.875 1.395 ;
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 1.275 0.475 1.445 1.015 ;
        RECT 3.435 0.475 3.605 1.015 ;
        RECT 1.275 0.305 3.605 0.475 ;
  END
END OAI21D1_3

#--------EOF---------

MACRO OR2D1
  CLASS CORE ;
  FOREIGN OR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.080 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.965400 ;
    PORT
      LAYER li1 ;
        RECT 3.355 2.545 3.685 2.715 ;
        RECT 3.435 1.185 3.605 2.545 ;
        RECT 3.355 1.015 3.685 1.185 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.735 2.275 2.065 2.445 ;
        RECT 1.815 1.765 1.985 2.275 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 0.000 -0.085 4.080 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 4.080 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 4.080 4.165 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 2.275 2.885 2.605 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 4.080 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 4.260 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.545 3.795 1.395 ;
      LAYER li1 ;
        RECT 0.115 2.545 3.065 2.715 ;
        RECT 2.895 2.445 3.065 2.545 ;
        RECT 2.815 2.275 3.145 2.445 ;
        RECT 1.195 1.935 1.525 2.105 ;
        RECT 1.275 1.185 1.445 1.935 ;
        RECT 2.895 1.765 3.065 2.275 ;
        RECT 2.815 1.595 3.145 1.765 ;
        RECT 1.195 1.015 1.525 1.185 ;
  END
END OR2D1

#--------EOF---------

MACRO OR2D1_1
  CLASS CORE ;
  FOREIGN OR2D1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.969900 ;
    PORT
      LAYER li1 ;
        RECT 3.355 2.545 3.685 2.715 ;
        RECT 3.435 1.185 3.605 2.545 ;
        RECT 3.355 1.015 3.685 1.185 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 2.355 0.085 2.525 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 0.000 -0.085 5.440 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 5.440 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 5.440 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 5.620 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.545 4.875 1.395 ;
      LAYER li1 ;
        RECT 2.275 2.545 2.605 2.715 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 2.275 2.275 2.605 2.445 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 1.275 0.475 1.445 1.015 ;
        RECT 1.195 0.305 1.525 0.475 ;
  END
END OR2D1_1

#--------EOF---------

MACRO OR2D1_2
  CLASS CORE ;
  FOREIGN OR2D1_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.965400 ;
    PORT
      LAYER li1 ;
        RECT 2.815 2.885 3.685 3.055 ;
        RECT 2.815 1.015 3.685 1.185 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 2.105 0.905 2.445 ;
        RECT 0.655 1.935 0.985 2.105 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.105 1.985 2.445 ;
        RECT 1.735 1.935 2.065 2.105 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 0.000 -0.085 5.440 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 5.440 4.165 ;
        RECT 2.355 3.055 2.525 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 5.440 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 5.620 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.545 4.875 1.395 ;
      LAYER li1 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 0.195 1.765 0.365 2.545 ;
        RECT 3.895 2.275 4.225 2.445 ;
        RECT 3.975 1.765 4.145 2.275 ;
        RECT 0.195 1.595 4.145 1.765 ;
        RECT 0.195 1.185 0.365 1.595 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 0.195 0.475 0.365 1.015 ;
        RECT 0.115 0.305 0.445 0.475 ;
  END
END OR2D1_2

#--------EOF---------

MACRO OR2D1_3
  CLASS CORE ;
  FOREIGN OR2D1_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.440 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.965400 ;
    PORT
      LAYER li1 ;
        RECT 2.815 2.545 3.685 2.715 ;
        RECT 2.815 1.015 3.685 1.185 ;
    END
  END z
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 1.815 1.765 1.985 2.105 ;
        RECT 1.735 1.595 2.065 1.765 ;
    END
  END a1
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.238500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 0.000 -0.085 5.440 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 5.440 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 5.440 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 5.440 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 5.620 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.545 4.875 1.395 ;
      LAYER li1 ;
        RECT 2.275 2.545 2.605 2.715 ;
        RECT 2.355 2.445 2.525 2.545 ;
        RECT 2.355 2.275 4.225 2.445 ;
        RECT 2.355 1.185 2.525 2.275 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 0.195 0.475 0.365 1.015 ;
        RECT 2.355 0.475 2.525 1.015 ;
        RECT 0.115 0.305 0.445 0.475 ;
        RECT 2.275 0.305 2.605 0.475 ;
  END
END OR2D1_3

#--------EOF---------

MACRO TIEH
  CLASS CORE ;
  FOREIGN TIEH ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.040 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.195 2.545 0.365 3.775 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 0.000 -0.085 2.040 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 2.040 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 2.040 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 2.040 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 2.220 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 1.635 1.395 ;
      LAYER li1 ;
        RECT 0.655 1.595 0.985 1.765 ;
        RECT 0.735 1.185 0.905 1.595 ;
        RECT 0.115 1.015 0.905 1.185 ;
  END
END TIEH

#--------EOF---------

MACRO TIEL
  CLASS CORE ;
  FOREIGN TIEL ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.040 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.195 1.015 0.905 1.185 ;
        RECT 0.735 0.305 0.905 1.015 ;
    END
  END zn
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 1.275 0.085 1.445 1.015 ;
        RECT 0.000 -0.085 2.040 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 2.040 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 2.040 4.165 ;
        RECT 1.275 3.055 1.445 3.995 ;
        RECT 1.195 2.885 1.525 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 2.040 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 2.220 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.485 1.635 1.395 ;
      LAYER li1 ;
        RECT 0.115 2.545 0.445 2.715 ;
        RECT 0.195 1.765 0.365 2.545 ;
        RECT 0.195 1.595 0.985 1.765 ;
  END
END TIEL

#--------EOF---------

MACRO XNR2D1
  CLASS CORE ;
  FOREIGN XNR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.735 1.765 0.905 2.105 ;
        RECT 0.655 1.595 0.985 1.765 ;
    END
  END a2
  PIN zn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 6.595 2.545 6.925 2.715 ;
        RECT 6.675 1.185 6.845 2.545 ;
        RECT 6.595 1.015 6.925 1.185 ;
    END
  END zn
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.276000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 2.545 2.605 2.715 ;
        RECT 2.355 1.765 2.525 2.545 ;
        RECT 1.735 1.595 2.525 1.765 ;
    END
  END a1
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 0.000 -0.085 8.500 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.500 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 8.500 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 8.500 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 8.680 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 8.115 1.395 ;
        RECT 0.005 0.485 1.635 0.715 ;
        RECT 6.485 0.485 8.115 0.715 ;
      LAYER li1 ;
        RECT 1.275 3.605 4.145 3.775 ;
        RECT 1.275 3.055 1.445 3.605 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 3.975 2.715 4.145 3.605 ;
        RECT 1.195 2.545 1.525 2.715 ;
        RECT 3.895 2.545 4.225 2.715 ;
        RECT 1.275 1.185 1.445 2.545 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 3.435 2.715 3.605 2.885 ;
        RECT 3.355 2.545 3.685 2.715 ;
        RECT 3.355 1.595 3.685 1.765 ;
        RECT 3.435 1.185 3.605 1.595 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 2.275 2.885 3.065 3.055 ;
        RECT 2.895 2.445 3.065 2.885 ;
        RECT 2.895 2.275 5.845 2.445 ;
        RECT 2.895 1.185 3.065 2.275 ;
        RECT 2.275 1.015 3.065 1.185 ;
        RECT 5.515 3.605 5.845 3.775 ;
        RECT 5.595 3.055 5.765 3.605 ;
        RECT 5.515 2.885 6.305 3.055 ;
        RECT 6.135 1.185 6.305 2.885 ;
        RECT 5.515 1.015 6.305 1.185 ;
  END
END XNR2D1

#--------EOF---------

MACRO XOR2D1
  CLASS CORE ;
  FOREIGN XOR2D1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.500 BY 4.080 ;
  SYMMETRY X Y R90 ;
  SITE obssite ;
  PIN a1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.291500 ;
    PORT
      LAYER li1 ;
        RECT 2.815 2.275 4.765 2.445 ;
        RECT 2.895 2.105 3.065 2.275 ;
        RECT 1.735 1.935 4.765 2.105 ;
    END
  END a1
  PIN z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006500 ;
    PORT
      LAYER li1 ;
        RECT 6.595 2.545 6.925 2.715 ;
        RECT 6.675 1.185 6.845 2.545 ;
        RECT 6.595 1.015 6.925 1.185 ;
    END
  END z
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.015 0.445 1.185 ;
        RECT 4.435 1.015 4.765 1.185 ;
        RECT 7.675 1.015 8.005 1.185 ;
        RECT 0.195 0.085 0.365 1.015 ;
        RECT 4.515 0.085 4.685 1.015 ;
        RECT 7.755 0.085 7.925 1.015 ;
        RECT 0.000 -0.085 8.500 0.085 ;
      LAYER mcon ;
        RECT 0.085 -0.085 0.255 0.085 ;
        RECT 0.425 -0.085 0.595 0.085 ;
        RECT 0.765 -0.085 0.935 0.085 ;
        RECT 1.105 -0.085 1.275 0.085 ;
        RECT 1.445 -0.085 1.615 0.085 ;
        RECT 1.785 -0.085 1.955 0.085 ;
        RECT 2.125 -0.085 2.295 0.085 ;
        RECT 2.465 -0.085 2.635 0.085 ;
        RECT 2.805 -0.085 2.975 0.085 ;
        RECT 3.145 -0.085 3.315 0.085 ;
        RECT 3.485 -0.085 3.655 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.165 -0.085 4.335 0.085 ;
        RECT 4.505 -0.085 4.675 0.085 ;
        RECT 4.845 -0.085 5.015 0.085 ;
        RECT 5.185 -0.085 5.355 0.085 ;
        RECT 5.525 -0.085 5.695 0.085 ;
        RECT 5.865 -0.085 6.035 0.085 ;
        RECT 6.205 -0.085 6.375 0.085 ;
        RECT 6.545 -0.085 6.715 0.085 ;
        RECT 6.885 -0.085 7.055 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
        RECT 7.565 -0.085 7.735 0.085 ;
        RECT 7.905 -0.085 8.075 0.085 ;
        RECT 8.245 -0.085 8.415 0.085 ;
      LAYER met1 ;
        RECT 0.000 -0.135 8.500 0.135 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 3.995 8.500 4.165 ;
        RECT 0.195 3.055 0.365 3.995 ;
        RECT 4.515 3.055 4.685 3.995 ;
        RECT 7.755 3.055 7.925 3.995 ;
        RECT 0.115 2.885 0.445 3.055 ;
        RECT 4.435 2.885 4.765 3.055 ;
        RECT 7.675 2.885 8.005 3.055 ;
      LAYER mcon ;
        RECT 0.085 3.995 0.255 4.165 ;
        RECT 0.425 3.995 0.595 4.165 ;
        RECT 0.765 3.995 0.935 4.165 ;
        RECT 1.105 3.995 1.275 4.165 ;
        RECT 1.445 3.995 1.615 4.165 ;
        RECT 1.785 3.995 1.955 4.165 ;
        RECT 2.125 3.995 2.295 4.165 ;
        RECT 2.465 3.995 2.635 4.165 ;
        RECT 2.805 3.995 2.975 4.165 ;
        RECT 3.145 3.995 3.315 4.165 ;
        RECT 3.485 3.995 3.655 4.165 ;
        RECT 3.825 3.995 3.995 4.165 ;
        RECT 4.165 3.995 4.335 4.165 ;
        RECT 4.505 3.995 4.675 4.165 ;
        RECT 4.845 3.995 5.015 4.165 ;
        RECT 5.185 3.995 5.355 4.165 ;
        RECT 5.525 3.995 5.695 4.165 ;
        RECT 5.865 3.995 6.035 4.165 ;
        RECT 6.205 3.995 6.375 4.165 ;
        RECT 6.545 3.995 6.715 4.165 ;
        RECT 6.885 3.995 7.055 4.165 ;
        RECT 7.225 3.995 7.395 4.165 ;
        RECT 7.565 3.995 7.735 4.165 ;
        RECT 7.905 3.995 8.075 4.165 ;
        RECT 8.245 3.995 8.415 4.165 ;
      LAYER met1 ;
        RECT 0.000 3.945 8.500 4.215 ;
    END
  END vdd
  OBS
      LAYER nwell ;
        RECT -0.180 1.865 8.680 4.405 ;
      LAYER pwell ;
        RECT 0.005 0.715 8.115 1.395 ;
        RECT 3.245 0.485 4.875 0.715 ;
        RECT 6.485 0.485 8.115 0.715 ;
      LAYER li1 ;
        RECT 1.195 2.885 1.525 3.055 ;
        RECT 1.275 1.185 1.445 2.885 ;
        RECT 1.195 1.015 1.525 1.185 ;
        RECT 2.275 3.605 2.605 3.775 ;
        RECT 4.975 3.605 7.465 3.775 ;
        RECT 2.355 3.055 2.525 3.605 ;
        RECT 2.275 2.885 2.605 3.055 ;
        RECT 5.055 1.765 5.225 3.605 ;
        RECT 2.355 1.595 5.225 1.765 ;
        RECT 2.355 1.185 2.525 1.595 ;
        RECT 2.275 1.015 2.605 1.185 ;
        RECT 1.735 3.605 2.065 3.775 ;
        RECT 1.815 2.715 1.985 3.605 ;
        RECT 3.355 2.885 3.685 3.055 ;
        RECT 3.435 2.715 3.605 2.885 ;
        RECT 1.815 2.545 3.605 2.715 ;
        RECT 3.355 1.015 3.685 1.185 ;
        RECT 3.435 0.475 3.605 1.015 ;
        RECT 0.655 0.305 3.605 0.475 ;
        RECT 5.515 2.885 5.845 3.055 ;
        RECT 5.595 1.185 5.765 2.885 ;
        RECT 5.515 1.015 5.845 1.185 ;
        RECT 5.595 0.475 5.765 1.015 ;
        RECT 5.515 0.305 5.845 0.475 ;
  END
END XOR2D1

#--------EOF---------


END LIBRARY
